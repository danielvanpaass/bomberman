library IEEE;
use IEEE.std_logic_1164.ALL;

entity tile_stdcrate_tb is
end tile_stdcrate_tb;

