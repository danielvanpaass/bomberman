library IEEE;
use IEEE.std_logic_1164.ALL;

entity hitbox_tb is
end hitbox_tb;

