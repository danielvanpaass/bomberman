configuration uneven_bits_behaviour_cfg of uneven_bits is
   for behaviour
   end for;
end uneven_bits_behaviour_cfg;
