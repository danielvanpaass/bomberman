configuration toplvl_coor_tb_behaviour_cfg of toplvl_coor_tb is
   for behaviour
      for all: toplvl_coor use configuration work.toplvl_coor_behaviour_cfg;
      end for;
   end for;
end toplvl_coor_tb_behaviour_cfg;
