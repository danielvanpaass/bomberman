configuration last_bomb_behaviour_cfg of last_bomb is
   for behaviour
   end for;
end last_bomb_behaviour_cfg;
