configuration toplvl_coor_behaviour_cfg of toplvl_coor is
   for behaviour
   end for;
end toplvl_coor_behaviour_cfg;
