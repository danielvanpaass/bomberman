library IEEE;
use IEEE.std_logic_1164.ALL;

architecture map_gen_behaviour of map_gen is
begin

end map_gen_behaviour;

