configuration selector_tb_behaviour_cfg of selector_tb is
   for behaviour
      for all: selector use configuration work.selector_behaviour_cfg;
      end for;
   end for;
end selector_tb_behaviour_cfg;
