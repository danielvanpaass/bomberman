configuration bombcook_behaviour_cfg of bombcook is
   for behaviour
   end for;
end bombcook_behaviour_cfg;
