library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour_bomb of hitbox_tb is
   component hitbox
      port(clk		 : in  std_logic;
   	reset	 : in  std_logic;
           crates   : in  std_logic_vector(120 downto 0);
           walls    : in  std_logic_vector(120 downto 0);
   	bomb_x_a	 : in  std_logic_vector(3 downto 0);
   	bomb_y_a	 : in  std_logic_vector(3 downto 0);
   	bomb_x_b	 : in  std_logic_vector(3 downto 0);
   	bomb_y_b	 : in  std_logic_vector(3 downto 0);
   	bomb_x_c	 : in  std_logic_vector(3 downto 0);
   	bomb_y_c	 : in  std_logic_vector(3 downto 0);
   	bomb_x_d	 : in  std_logic_vector(3 downto 0);
   	bomb_y_d	 : in  std_logic_vector(3 downto 0);
   	bomb_x_e	 : in  std_logic_vector(3 downto 0);
   	bomb_y_e	 : in  std_logic_vector(3 downto 0);
   	bomb_x_f	 : in  std_logic_vector(3 downto 0);
   	bomb_y_f	 : in  std_logic_vector(3 downto 0);
   	bomb_x_g	 : in  std_logic_vector(3 downto 0);
   	bomb_y_g	 : in  std_logic_vector(3 downto 0);
   	bomb_x_h	 : in  std_logic_vector(3 downto 0);
   	bomb_y_h	 : in  std_logic_vector(3 downto 0);
   	bomb_a_active : in std_logic;
   	bomb_b_active : in std_logic;
   	bomb_c_active : in std_logic;
   	bomb_d_active : in std_logic;
   	bomb_e_active : in std_logic;
   	bomb_f_active : in std_logic;
   	bomb_g_active : in std_logic;
   	bomb_h_active : in std_logic;
           right_p1 : in  std_logic;
           x_p1 : out std_logic_vector(3 downto 0);
           y_p1 : out std_logic_vector(3 downto 0));
   end component;
   signal clk		 : std_logic;
   signal reset	 : std_logic;
   signal crates   : std_logic_vector(120 downto 0);
   signal walls    : std_logic_vector(120 downto 0);
   signal bomb_x_a	 : std_logic_vector(3 downto 0);
   signal bomb_y_a	 : std_logic_vector(3 downto 0);
   signal bomb_x_b	 : std_logic_vector(3 downto 0);
   signal bomb_y_b	 : std_logic_vector(3 downto 0);
   signal bomb_x_c	 : std_logic_vector(3 downto 0);
   signal bomb_y_c	 : std_logic_vector(3 downto 0);
   signal bomb_x_d	 : std_logic_vector(3 downto 0);
   signal bomb_y_d	 : std_logic_vector(3 downto 0);
   signal bomb_x_e	 : std_logic_vector(3 downto 0);
   signal bomb_y_e	 : std_logic_vector(3 downto 0);
   signal bomb_x_f	 : std_logic_vector(3 downto 0);
   signal bomb_y_f	 : std_logic_vector(3 downto 0);
   signal bomb_x_g	 : std_logic_vector(3 downto 0);
   signal bomb_y_g	 : std_logic_vector(3 downto 0);
   signal bomb_x_h	 : std_logic_vector(3 downto 0);
   signal bomb_y_h	 : std_logic_vector(3 downto 0);
   signal bomb_a_active : std_logic;
   signal bomb_b_active : std_logic;
   signal bomb_c_active : std_logic;
   signal bomb_d_active : std_logic;
   signal bomb_e_active : std_logic;
   signal bomb_f_active : std_logic;
   signal bomb_g_active : std_logic;
   signal bomb_h_active : std_logic;
   signal right_p1 : std_logic;
   signal x_p1 : std_logic_vector(3 downto 0);
   signal y_p1 : std_logic_vector(3 downto 0);
begin
test: hitbox port map (clk, reset, crates, walls, bomb_x_a, bomb_y_a, bomb_x_b, bomb_y_b, bomb_x_c, bomb_y_c, bomb_x_d, bomb_y_d, bomb_x_e, bomb_y_e, bomb_x_f, bomb_y_f, bomb_x_g, bomb_y_g, bomb_x_h, bomb_y_h, bomb_a_active, bomb_b_active, bomb_c_active, bomb_d_active, bomb_e_active, bomb_f_active, bomb_g_active, bomb_h_active, right_p1, x_p1, y_p1);
clk <= '1' after 0 ns,
     '0' after 0.04 ms when clk /= '0' else '1' after 0.04 ms;

      reset <= '1' after 0 ns,
	 '0' after 0.12 ms;
   crates(0) <= '0' after 0 ns;
   crates(1) <= '0' after 0 ns;
   crates(2) <= '0' after 0 ns;
   crates(3) <= '0' after 0 ns;
   crates(4) <= '0' after 0 ns;
   crates(5) <= '0' after 0 ns;
   crates(6) <= '0' after 0 ns;
   crates(7) <= '0' after 0 ns;
   crates(8) <= '0' after 0 ns;
   crates(9) <= '0' after 0 ns;
   crates(10) <= '0' after 0 ns;
   crates(11) <= '0' after 0 ns;
   crates(12) <= '0' after 0 ns;
   crates(13) <= '0' after 0 ns;
   crates(14) <= '0' after 0 ns;
   crates(15) <= '0' after 0 ns;
   crates(16) <= '0' after 0 ns;
   crates(17) <= '0' after 0 ns;
   crates(18) <= '0' after 0 ns;
   crates(19) <= '0' after 0 ns;
   crates(20) <= '0' after 0 ns;
   crates(21) <= '0' after 0 ns;
   crates(22) <= '0' after 0 ns;
   crates(23) <= '0' after 0 ns;
   crates(24) <= '0' after 0 ns;
   crates(25) <= '0' after 0 ns;
   crates(26) <= '0' after 0 ns;
   crates(27) <= '0' after 0 ns;
   crates(28) <= '0' after 0 ns;
   crates(29) <= '0' after 0 ns;
   crates(30) <= '0' after 0 ns;
   crates(31) <= '0' after 0 ns;
   crates(32) <= '0' after 0 ns;
   crates(33) <= '0' after 0 ns;
   crates(34) <= '0' after 0 ns;
   crates(35) <= '0' after 0 ns;
   crates(36) <= '0' after 0 ns;
   crates(37) <= '0' after 0 ns;
   crates(38) <= '0' after 0 ns;
   crates(39) <= '0' after 0 ns;
   crates(40) <= '0' after 0 ns;
   crates(41) <= '0' after 0 ns;
   crates(42) <= '0' after 0 ns;
   crates(43) <= '0' after 0 ns;
   crates(44) <= '0' after 0 ns;
   crates(45) <= '0' after 0 ns;
   crates(46) <= '0' after 0 ns;
   crates(47) <= '0' after 0 ns;
   crates(48) <= '0' after 0 ns;
   crates(49) <= '0' after 0 ns;
   crates(50) <= '0' after 0 ns;
   crates(51) <= '0' after 0 ns;
   crates(52) <= '0' after 0 ns;
   crates(53) <= '0' after 0 ns;
   crates(54) <= '0' after 0 ns;
   crates(55) <= '0' after 0 ns;
   crates(56) <= '0' after 0 ns;
   crates(57) <= '0' after 0 ns;
   crates(58) <= '0' after 0 ns;
   crates(59) <= '0' after 0 ns;
   crates(60) <= '0' after 0 ns;
   crates(61) <= '0' after 0 ns;
   crates(62) <= '0' after 0 ns;
   crates(63) <= '0' after 0 ns;
   crates(64) <= '0' after 0 ns;
   crates(65) <= '0' after 0 ns;
   crates(66) <= '0' after 0 ns;
   crates(67) <= '0' after 0 ns;
   crates(68) <= '0' after 0 ns;
   crates(69) <= '0' after 0 ns;
   crates(70) <= '0' after 0 ns;
   crates(71) <= '0' after 0 ns;
   crates(72) <= '0' after 0 ns;
   crates(73) <= '0' after 0 ns;
   crates(74) <= '0' after 0 ns;
   crates(75) <= '0' after 0 ns;
   crates(76) <= '0' after 0 ns;
   crates(77) <= '0' after 0 ns;
   crates(78) <= '0' after 0 ns;
   crates(79) <= '0' after 0 ns;
   crates(80) <= '0' after 0 ns;
   crates(81) <= '0' after 0 ns;
   crates(82) <= '0' after 0 ns;
   crates(83) <= '0' after 0 ns;
   crates(84) <= '0' after 0 ns;
   crates(85) <= '0' after 0 ns;
   crates(86) <= '0' after 0 ns;
   crates(87) <= '0' after 0 ns;
   crates(88) <= '0' after 0 ns;
   crates(89) <= '0' after 0 ns;
   crates(90) <= '0' after 0 ns;
   crates(91) <= '0' after 0 ns;
   crates(92) <= '0' after 0 ns;
   crates(93) <= '0' after 0 ns;
   crates(94) <= '0' after 0 ns;
   crates(95) <= '0' after 0 ns;
   crates(96) <= '0' after 0 ns;
   crates(97) <= '0' after 0 ns;
   crates(98) <= '0' after 0 ns;
   crates(99) <= '0' after 0 ns;
   crates(100) <= '0' after 0 ns;
   crates(101) <= '0' after 0 ns;
   crates(102) <= '0' after 0 ns;
   crates(103) <= '0' after 0 ns;
   crates(104) <= '0' after 0 ns;
   crates(105) <= '0' after 0 ns;
   crates(106) <= '0' after 0 ns;
   crates(107) <= '0' after 0 ns;
   crates(108) <= '0' after 0 ns;
   crates(109) <= '0' after 0 ns;
   crates(110) <= '0' after 0 ns;
   crates(111) <= '0' after 0 ns;
   crates(112) <= '0' after 0 ns;
   crates(113) <= '0' after 0 ns;
   crates(114) <= '0' after 0 ns;
   crates(115) <= '0' after 0 ns;
   crates(116) <= '0' after 0 ns;
   crates(117) <= '0' after 0 ns;
   crates(118) <= '0' after 0 ns;
   crates(119) <= '0' after 0 ns;
   crates(120) <= '0' after 0 ns;
   walls(0) <= '0' after 0 ns;
   walls(1) <= '0' after 0 ns;
   walls(2) <= '0' after 0 ns;
   walls(3) <= '0' after 0 ns;
   walls(4) <= '0' after 0 ns;
   walls(5) <= '0' after 0 ns;
   walls(6) <= '0' after 0 ns;
   walls(7) <= '0' after 0 ns;
   walls(8) <= '0' after 0 ns;
   walls(9) <= '0' after 0 ns;
   walls(10) <= '0' after 0 ns;
   walls(11) <= '0' after 0 ns;
   walls(12) <= '0' after 0 ns;
   walls(13) <= '0' after 0 ns;
   walls(14) <= '0' after 0 ns;
   walls(15) <= '0' after 0 ns;
   walls(16) <= '0' after 0 ns;
   walls(17) <= '0' after 0 ns;
   walls(18) <= '0' after 0 ns;
   walls(19) <= '0' after 0 ns;
   walls(20) <= '0' after 0 ns;
   walls(21) <= '0' after 0 ns;
   walls(22) <= '0' after 0 ns;
   walls(23) <= '0' after 0 ns;
   walls(24) <= '0' after 0 ns;
   walls(25) <= '0' after 0 ns;
   walls(26) <= '0' after 0 ns;
   walls(27) <= '0' after 0 ns;
   walls(28) <= '0' after 0 ns;
   walls(29) <= '0' after 0 ns;
   walls(30) <= '0' after 0 ns;
   walls(31) <= '0' after 0 ns;
   walls(32) <= '0' after 0 ns;
   walls(33) <= '0' after 0 ns;
   walls(34) <= '0' after 0 ns;
   walls(35) <= '0' after 0 ns;
   walls(36) <= '0' after 0 ns;
   walls(37) <= '0' after 0 ns;
   walls(38) <= '0' after 0 ns;
   walls(39) <= '0' after 0 ns;
   walls(40) <= '0' after 0 ns;
   walls(41) <= '0' after 0 ns;
   walls(42) <= '0' after 0 ns;
   walls(43) <= '0' after 0 ns;
   walls(44) <= '0' after 0 ns;
   walls(45) <= '0' after 0 ns;
   walls(46) <= '0' after 0 ns;
   walls(47) <= '0' after 0 ns;
   walls(48) <= '0' after 0 ns;
   walls(49) <= '0' after 0 ns;
   walls(50) <= '0' after 0 ns;
   walls(51) <= '0' after 0 ns;
   walls(52) <= '0' after 0 ns;
   walls(53) <= '0' after 0 ns;
   walls(54) <= '0' after 0 ns;
   walls(55) <= '0' after 0 ns;
   walls(56) <= '0' after 0 ns;
   walls(57) <= '0' after 0 ns;
   walls(58) <= '0' after 0 ns;
   walls(59) <= '0' after 0 ns;
   walls(60) <= '0' after 0 ns;
   walls(61) <= '0' after 0 ns;
   walls(62) <= '0' after 0 ns;
   walls(63) <= '0' after 0 ns;
   walls(64) <= '0' after 0 ns;
   walls(65) <= '0' after 0 ns;
   walls(66) <= '0' after 0 ns;
   walls(67) <= '0' after 0 ns;
   walls(68) <= '0' after 0 ns;
   walls(69) <= '0' after 0 ns;
   walls(70) <= '0' after 0 ns;
   walls(71) <= '0' after 0 ns;
   walls(72) <= '0' after 0 ns;
   walls(73) <= '0' after 0 ns;
   walls(74) <= '0' after 0 ns;
   walls(75) <= '0' after 0 ns;
   walls(76) <= '0' after 0 ns;
   walls(77) <= '0' after 0 ns;
   walls(78) <= '0' after 0 ns;
   walls(79) <= '0' after 0 ns;
   walls(80) <= '0' after 0 ns;
   walls(81) <= '0' after 0 ns;
   walls(82) <= '0' after 0 ns;
   walls(83) <= '0' after 0 ns;
   walls(84) <= '0' after 0 ns;
   walls(85) <= '0' after 0 ns;
   walls(86) <= '0' after 0 ns;
   walls(87) <= '0' after 0 ns;
   walls(88) <= '0' after 0 ns;
   walls(89) <= '0' after 0 ns;
   walls(90) <= '0' after 0 ns;
   walls(91) <= '0' after 0 ns;
   walls(92) <= '0' after 0 ns;
   walls(93) <= '0' after 0 ns;
   walls(94) <= '0' after 0 ns;
   walls(95) <= '0' after 0 ns;
   walls(96) <= '0' after 0 ns;
   walls(97) <= '0' after 0 ns;
   walls(98) <= '0' after 0 ns;
   walls(99) <= '0' after 0 ns;
   walls(100) <= '0' after 0 ns;
   walls(101) <= '0' after 0 ns;
   walls(102) <= '0' after 0 ns;
   walls(103) <= '0' after 0 ns;
   walls(104) <= '0' after 0 ns;
   walls(105) <= '0' after 0 ns;
   walls(106) <= '0' after 0 ns;
   walls(107) <= '0' after 0 ns;
   walls(108) <= '0' after 0 ns;
   walls(109) <= '0' after 0 ns;
   walls(110) <= '0' after 0 ns;
   walls(111) <= '0' after 0 ns;
   walls(112) <= '0' after 0 ns;
   walls(113) <= '0' after 0 ns;
   walls(114) <= '0' after 0 ns;
   walls(115) <= '0' after 0 ns;
   walls(116) <= '0' after 0 ns;
   walls(117) <= '0' after 0 ns;
   walls(118) <= '0' after 0 ns;
   walls(119) <= '0' after 0 ns;
   walls(120) <= '0' after 0 ns;
   bomb_x_a(0) <= '0' after 0 ns;
   bomb_x_a(1) <= '0' after 0 ns;
   bomb_x_a(2) <= '1' after 0 ns;
   bomb_x_a(3) <= '0' after 0 ns;
   bomb_y_a(0) <= '0' after 0 ns;
   bomb_y_a(1) <= '0' after 0 ns;
   bomb_y_a(2) <= '0' after 0 ns;
   bomb_y_a(3) <= '0' after 0 ns;
   bomb_x_b(0) <= '0' after 0 ns;
   bomb_x_b(1) <= '0' after 0 ns;
   bomb_x_b(2) <= '0' after 0 ns;
   bomb_x_b(3) <= '0' after 0 ns;
   bomb_y_b(0) <= '0' after 0 ns;
   bomb_y_b(1) <= '0' after 0 ns;
   bomb_y_b(2) <= '0' after 0 ns;
   bomb_y_b(3) <= '0' after 0 ns;
   bomb_x_c(0) <= '0' after 0 ns;
   bomb_x_c(1) <= '0' after 0 ns;
   bomb_x_c(2) <= '0' after 0 ns;
   bomb_x_c(3) <= '0' after 0 ns;
   bomb_y_c(0) <= '0' after 0 ns;
   bomb_y_c(1) <= '0' after 0 ns;
   bomb_y_c(2) <= '0' after 0 ns;
   bomb_y_c(3) <= '0' after 0 ns;
   bomb_x_d(0) <= '0' after 0 ns;
   bomb_x_d(1) <= '0' after 0 ns;
   bomb_x_d(2) <= '0' after 0 ns;
   bomb_x_d(3) <= '0' after 0 ns;
   bomb_y_d(0) <= '0' after 0 ns;
   bomb_y_d(1) <= '0' after 0 ns;
   bomb_y_d(2) <= '0' after 0 ns;
   bomb_y_d(3) <= '0' after 0 ns;
   bomb_x_e(0) <= '0' after 0 ns;
   bomb_x_e(1) <= '0' after 0 ns;
   bomb_x_e(2) <= '0' after 0 ns;
   bomb_x_e(3) <= '0' after 0 ns;
   bomb_y_e(0) <= '0' after 0 ns;
   bomb_y_e(1) <= '0' after 0 ns;
   bomb_y_e(2) <= '0' after 0 ns;
   bomb_y_e(3) <= '0' after 0 ns;
   bomb_x_f(0) <= '0' after 0 ns;
   bomb_x_f(1) <= '0' after 0 ns;
   bomb_x_f(2) <= '0' after 0 ns;
   bomb_x_f(3) <= '0' after 0 ns;
   bomb_y_f(0) <= '0' after 0 ns;
   bomb_y_f(1) <= '0' after 0 ns;
   bomb_y_f(2) <= '0' after 0 ns;
   bomb_y_f(3) <= '0' after 0 ns;
   bomb_x_g(0) <= '0' after 0 ns;
   bomb_x_g(1) <= '0' after 0 ns;
   bomb_x_g(2) <= '0' after 0 ns;
   bomb_x_g(3) <= '0' after 0 ns;
   bomb_y_g(0) <= '0' after 0 ns;
   bomb_y_g(1) <= '0' after 0 ns;
   bomb_y_g(2) <= '0' after 0 ns;
   bomb_y_g(3) <= '0' after 0 ns;
   bomb_x_h(0) <= '0' after 0 ns;
   bomb_x_h(1) <= '0' after 0 ns;
   bomb_x_h(2) <= '0' after 0 ns;
   bomb_x_h(3) <= '0' after 0 ns;
   bomb_y_h(0) <= '0' after 0 ns;
   bomb_y_h(1) <= '0' after 0 ns;
   bomb_y_h(2) <= '0' after 0 ns;
   bomb_y_h(3) <= '0' after 0 ns;
   bomb_a_active <= '0' after 0 ns,
   '1' after 250 ms;
   bomb_b_active <= '0' after 0 ns;
   bomb_c_active <= '0' after 0 ns;
   bomb_d_active <= '0' after 0 ns;
   bomb_e_active <= '0' after 0 ns;
   bomb_f_active <= '0' after 0 ns;
   bomb_g_active <= '0' after 0 ns;
   bomb_h_active <= '0' after 0 ns;
 right_p1 <= '0' after 0 ns,
		'1' after 100 ns,
'0' after 200 ns,
'1' after 800 ns,
'0' after 1400 ns,
'1' after 1800 ns;

end behaviour_bomb;

