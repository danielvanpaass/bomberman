library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of playground is

component tile_stdempty is
   port(xlethal : in  std_logic;
	ylethal : in std_logic;
	expl : in std_logic;
	clk : in std_logic;
	reset : in std_logic;
	tiletype : out std_logic_vector(1 downto 0));
end component;

component tile_stdcrate is
   port(xlethal : in  std_logic;
	ylethal : in std_logic;
	expl : in std_logic;
	clk : in std_logic;
	reset : in std_logic;
	tiletype : out std_logic_vector(1 downto 0));
end component;

component xy_convert is
   port(x_in : in  std_logic_vector(3 downto 0);
	y_in : in  std_logic_vector(3 downto 0);
	x0 : out std_logic;
	x1 : out std_logic;
	x2 : out std_logic;
	x3 : out std_logic;
	x4 : out std_logic;
	x5 : out std_logic;
	x6 : out std_logic;
	x7 : out std_logic;
	x8 : out std_logic;
	x9 : out std_logic;
	x10 : out std_logic;
	y0 : out std_logic;
	y1 : out std_logic;
	y2 : out std_logic;
	y3 : out std_logic;
	y4 : out std_logic;
	y5 : out std_logic;
	y6 : out std_logic;
	y7 : out std_logic;
	y8 : out std_logic;
	y9 : out std_logic;
	y10 : out std_logic);
end component;

signal xo0, xo1, xo2, xo3, xo4, xo5, xo6, xo7, xo8, xo9,xo10,yo0, yo1, yo2, yo3, yo4, yo5, yo6, yo7, yo8, yo9,yo10: std_logic;

begin
--xy conversion to call seperate fsms
xyconv: xy_convert port map(lethalx, lethaly,xo0, xo1, xo2, xo3, xo4, xo5, xo6, xo7, xo8, xo9,xo10,yo0, yo1, yo2, yo3, yo4, yo5, yo6, yo7, yo8, yo9,yo10);

--this was made to solve a warning with quartus
xo0<='1';
xo10<='1';
yo0<='1';
yo10<='1';

--t1 to t11, for y1, "1111111111111111111111", all walls
t1to11: y0 <= "1111111111111111111111";

--t12 to t22, t12 and t22 being "00" (walls)
y1(21) <= '1'; --t12
y1(20) <= '1';
t13: tile_stdempty port map(xo1, yo1, lethal, clk, reset => reset, tiletype(1) => y1(19), tiletype(0) => y1(18));
t14: tile_stdempty port map(xo2, yo1, lethal, clk, reset => reset, tiletype(1) => y1(17), tiletype(0) => y1(16));
t15: tile_stdempty port map(xo3, yo1, lethal, clk, reset => reset, tiletype(1) => y1(15), tiletype(0) => y1(14));
t16: tile_stdcrate port map(xo4, yo1, lethal, clk, reset => reset, tiletype(1) => y1(13), tiletype(0) => y1(12));
t17: tile_stdcrate port map(xo5, yo1, lethal, clk, reset => reset, tiletype(1) => y1(11), tiletype(0) => y1(10));
t18: tile_stdcrate port map(xo6, yo1, lethal, clk, reset => reset, tiletype(1) => y1(9), tiletype(0) => y1(8));
t19: tile_stdempty port map(xo7, yo1, lethal, clk, reset => reset, tiletype(1) => y1(7), tiletype(0) => y1(6));
t20: tile_stdempty port map(xo8, yo1, lethal, clk, reset => reset, tiletype(1) => y1(5), tiletype(0) => y1(4));
t21: tile_stdempty port map(xo9, yo1, lethal, clk, reset => reset, tiletype(1) => y1(3), tiletype(0) => y1(2));
y1(1) <= '1'; --t22
y1(0) <= '1';

--t23 to t33, t23 and t33 being "00" (walls)
y2(21) <= '1'; --t23
y2(20) <= '1';
t24: tile_stdempty port map(xo1, yo2, lethal, clk, reset => reset, tiletype(1) => y2(19), tiletype(0) => y2(18));
y2(17) <= '1'; --wall
y2(16) <= '1'; --wall
t26: tile_stdcrate port map(xo3, yo2, lethal, clk, reset => reset, tiletype(1) => y2(15), tiletype(0) => y2(14));
y2(13) <= '1'; --wall
y2(12) <= '1'; --wall
t28: tile_stdcrate port map(xo5, yo2, lethal, clk, reset => reset, tiletype(1) => y2(11), tiletype(0) => y2(10));
y2(9) <= '1'; --wall
y2(8) <= '1'; --wall
t30: tile_stdcrate port map(xo7, yo2, lethal, clk, reset => reset, tiletype(1) => y2(7), tiletype(0) => y2(6));
y2(5) <= '1'; --wall
y2(4) <= '1'; --wall
t32: tile_stdempty port map(xo9, yo2, lethal, clk, reset => reset, tiletype(1) => y2(3), tiletype(0) => y2(2));
y2(1) <= '1'; --t33
y2(0) <= '1';

--t34 to t44
y3(21) <= '1'; --wall
y3(20) <= '1'; --wall
t35: tile_stdempty port map(xo1, yo3, lethal, clk, reset => reset, tiletype(1) => y3(19), tiletype(0) => y3(18));
t36: tile_stdcrate port map(xo2, yo3, lethal, clk, reset => reset, tiletype(1) => y3(17), tiletype(0) => y3(16));
t37: tile_stdcrate port map(xo3, yo3, lethal, clk, reset => reset, tiletype(1) => y3(15), tiletype(0) => y3(14));
t38: tile_stdcrate port map(xo4, yo3, lethal, clk, reset => reset, tiletype(1) => y3(13), tiletype(0) => y3(12));
t39: tile_stdcrate port map(xo5, yo3, lethal, clk, reset => reset, tiletype(1) => y3(11), tiletype(0) => y3(10));
t40: tile_stdcrate port map(xo6, yo3, lethal, clk, reset => reset, tiletype(1) => y3(9), tiletype(0) => y3(8));
t41: tile_stdcrate port map(xo7, yo3, lethal, clk, reset => reset, tiletype(1) => y3(7), tiletype(0) => y3(6));
t42: tile_stdcrate port map(xo8, yo3, lethal, clk, reset => reset, tiletype(1) => y3(5), tiletype(0) => y3(4));
t43: tile_stdempty port map(xo9, yo3, lethal, clk, reset => reset, tiletype(1) => y3(3), tiletype(0) => y3(2));
y3(1) <= '1'; --wall
y3(0) <= '1'; --wall

--t45 to t55
y4(21) <= '1'; 
y4(20) <= '1';
t46: tile_stdcrate port map(xo1, yo4, lethal, clk, reset => reset, tiletype(1) => y4(19), tiletype(0) => y4(18));
y4(17) <= '1'; --wall
y4(16) <= '1'; --wall
t48: tile_stdcrate port map(xo3, yo4, lethal, clk, reset => reset, tiletype(1) => y4(15), tiletype(0) => y4(14));
y4(13) <= '1'; --wall
y4(12) <= '1'; --wall
t50: tile_stdempty port map(xo5, yo4, lethal, clk, reset => reset, tiletype(1) => y4(11), tiletype(0) => y4(10));
y4(9) <= '1'; --wall
y4(8) <= '1'; --wall
t52: tile_stdcrate port map(xo7, yo4, lethal, clk, reset => reset, tiletype(1) => y4(7), tiletype(0) => y4(6));
y4(5) <= '1'; --wall
y4(4) <= '1'; --wall
t54: tile_stdcrate port map(xo9, yo4, lethal, clk, reset => reset, tiletype(1) => y4(3), tiletype(0) => y4(2));
y4(1) <= '1'; 
y4(0) <= '1';

--t56 to t66
y5(21) <= '1'; --wall
y5(20) <= '1'; --wall
t57: tile_stdcrate port map(xo1, yo5, lethal, clk, reset => reset, tiletype(1) => y5(19), tiletype(0) => y5(18));
t58: tile_stdcrate port map(xo2, yo5, lethal, clk, reset => reset, tiletype(1) => y5(17), tiletype(0) => y5(16));
t59: tile_stdcrate port map(xo3, yo5, lethal, clk, reset => reset, tiletype(1) => y5(15), tiletype(0) => y5(14));
t60: tile_stdempty port map(xo4, yo5, lethal, clk, reset => reset, tiletype(1) => y5(13), tiletype(0) => y5(12));
t61: tile_stdempty port map(xo5, yo5, lethal, clk, reset => reset, tiletype(1) => y5(11), tiletype(0) => y5(10));
t62: tile_stdempty port map(xo6, yo5, lethal, clk, reset => reset, tiletype(1) => y5(9), tiletype(0) => y5(8));
t63: tile_stdcrate port map(xo7, yo5, lethal, clk, reset => reset, tiletype(1) => y5(7), tiletype(0) => y5(6));
t64: tile_stdcrate port map(xo8, yo5, lethal, clk, reset => reset, tiletype(1) => y5(5), tiletype(0) => y5(4));
t65: tile_stdcrate port map(xo9, yo5, lethal, clk, reset => reset, tiletype(1) => y5(3), tiletype(0) => y5(2));
y5(1) <= '1'; --wall
y5(0) <= '1'; --wall

--t67 to t77
y6(21) <= '1'; 
y6(20) <= '1';
t68: tile_stdcrate port map(xo1, yo6, lethal, clk, reset => reset, tiletype(1) => y6(19), tiletype(0) => y6(18));
y6(17) <= '1'; --wall
y6(16) <= '1'; --wall
t70: tile_stdcrate port map(xo3, yo6, lethal, clk, reset => reset, tiletype(1) => y6(15), tiletype(0) => y6(14));
y6(13) <= '1'; --wall
y6(12) <= '1'; --wall
t72: tile_stdempty port map(xo5, yo6, lethal, clk, reset => reset, tiletype(1) => y6(11), tiletype(0) => y6(10));
y6(9) <= '1'; --wall
y6(8) <= '1'; --wall
t74: tile_stdcrate port map(xo7, yo6, lethal, clk, reset => reset, tiletype(1) => y6(7), tiletype(0) => y6(6));
y6(5) <= '1'; --wall
y6(4) <= '1'; --wall
t76: tile_stdcrate port map(xo9, yo6, lethal, clk, reset => reset, tiletype(1) => y6(3), tiletype(0) => y6(2));
y6(1) <= '1'; 
y6(0) <= '1';

--t78 to t88
y7(21) <= '1'; --wall
y7(20) <= '1'; --wall
t79: tile_stdempty port map(xo1, yo7, lethal, clk, reset => reset, tiletype(1) => y7(19), tiletype(0) => y7(18));
t80: tile_stdcrate port map(xo2, yo7, lethal, clk, reset => reset, tiletype(1) => y7(17), tiletype(0) => y7(16));
t81: tile_stdcrate port map(xo3, yo7, lethal, clk, reset => reset, tiletype(1) => y7(15), tiletype(0) => y7(14));
t82: tile_stdcrate port map(xo4, yo7, lethal, clk, reset => reset, tiletype(1) => y7(13), tiletype(0) => y7(12));
t83: tile_stdcrate port map(xo5, yo7, lethal, clk, reset => reset, tiletype(1) => y7(11), tiletype(0) => y7(10));
t84: tile_stdcrate port map(xo6, yo7, lethal, clk, reset => reset, tiletype(1) => y7(9), tiletype(0) => y7(8));
t85: tile_stdcrate port map(xo7, yo7, lethal, clk, reset => reset, tiletype(1) => y7(7), tiletype(0) => y7(6));
t86: tile_stdcrate port map(xo8, yo7, lethal, clk, reset => reset, tiletype(1) => y7(5), tiletype(0) => y7(4));
t87: tile_stdempty port map(xo9, yo7, lethal, clk, reset => reset, tiletype(1) => y7(3), tiletype(0) => y7(2));
y7(1) <= '1'; --wall
y7(0) <= '1'; --wall

--t89 to t99
y8(21) <= '1';
y8(20) <= '1';
t90: tile_stdempty port map(xo1, yo8, lethal, clk, reset => reset, tiletype(1) => y8(19), tiletype(0) => y8(18));
y8(17) <= '1'; --wall
y8(16) <= '1'; --wall
t92: tile_stdcrate port map(xo3, yo8, lethal, clk, reset => reset, tiletype(1) => y8(15), tiletype(0) => y8(14));
y8(13) <= '1'; --wall
y8(12) <= '1'; --wall
t94: tile_stdcrate port map(xo5, yo8, lethal, clk, reset => reset, tiletype(1) => y8(11), tiletype(0) => y8(10));
y8(9) <= '1'; --wall
y8(8) <= '1'; --wall
t96: tile_stdcrate port map(xo7, yo8, lethal, clk, reset => reset, tiletype(1) => y8(7), tiletype(0) => y8(6));
y8(5) <= '1'; --wall
y8(4) <= '1'; --wall
t98: tile_stdempty port map(xo9, yo8, lethal, clk, reset => reset, tiletype(1) => y8(3), tiletype(0) => y8(2));
y8(1) <= '1'; --t33
y8(0) <= '1';

--t100 to t110
y9(21) <= '1';
y9(20) <= '1';
t101: tile_stdempty port map(xo1, yo9, lethal, clk, reset => reset, tiletype(1) => y9(19), tiletype(0) => y9(18));
t102: tile_stdempty port map(xo2, yo9, lethal, clk, reset => reset, tiletype(1) => y9(17), tiletype(0) => y9(16));
t103: tile_stdempty port map(xo3, yo9, lethal, clk, reset => reset, tiletype(1) => y9(15), tiletype(0) => y9(14));
t104: tile_stdcrate port map(xo4, yo9, lethal, clk, reset => reset, tiletype(1) => y9(13), tiletype(0) => y9(12));
t105: tile_stdcrate port map(xo5, yo9, lethal, clk, reset => reset, tiletype(1) => y9(11), tiletype(0) => y9(10));
t106: tile_stdcrate port map(xo6, yo9, lethal, clk, reset => reset, tiletype(1) => y9(9), tiletype(0) => y9(8));
t107: tile_stdempty port map(xo7, yo9, lethal, clk, reset => reset, tiletype(1) => y9(7), tiletype(0) => y9(6));
t108: tile_stdempty port map(xo8, yo9, lethal, clk, reset => reset, tiletype(1) => y9(5), tiletype(0) => y9(4));
t109: tile_stdempty port map(xo9, yo9, lethal, clk, reset => reset, tiletype(1) => y9(3), tiletype(0) => y9(2));
y9(1) <= '1';
y9(0) <= '1';

--t111 to t121, for y10, "1111111111111111111111", all walls
t111to121: y10 <= "1111111111111111111111";

end behaviour;

