
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of toplvl_coor is

  component BUFFD1P5BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component BUFFD2BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCNQD1BWP7T
    port(CP, CN, D : in std_logic; Q : out std_logic);
  end component;

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component MOAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component OAI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component INR2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component DFKCND1BWP7T
    port(CP, CN, D : in std_logic; Q, QN : out std_logic);
  end component;

  component AN2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component BUFFD4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component AN2D4BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component LHQD1BWP7T
    port(E, D : in std_logic; Q : out std_logic);
  end component;

  component AO221D0BWP7T
    port(A1, A2, B1, B2, C : in std_logic; Z : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component INVD4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component CKAN2D8BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component TIELBWP7T
    port(ZN : out std_logic);
  end component;

  component TIEHBWP7T
    port(Z : out std_logic);
  end component;

  signal bombnop1 : std_logic_vector(3 downto 0);
  signal bombselp1_state : std_logic_vector(2 downto 0);
  signal bombnop2 : std_logic_vector(3 downto 0);
  signal bombselp2_state : std_logic_vector(2 downto 0);
  signal bombcooka_state : std_logic_vector(1 downto 0);
  signal bombcooka_bombxsample : std_logic_vector(3 downto 0);
  signal bombcooka_bombysample : std_logic_vector(3 downto 0);
  signal bombcookb_state : std_logic_vector(1 downto 0);
  signal bombcookb_bombxsample : std_logic_vector(3 downto 0);
  signal bombcookb_bombysample : std_logic_vector(3 downto 0);
  signal bombcookc_state : std_logic_vector(1 downto 0);
  signal bombcookc_bombxsample : std_logic_vector(3 downto 0);
  signal bombcookc_bombysample : std_logic_vector(3 downto 0);
  signal bombcookd_state : std_logic_vector(1 downto 0);
  signal bombcookd_bombxsample : std_logic_vector(3 downto 0);
  signal bombcookd_bombysample : std_logic_vector(3 downto 0);
  signal bombcooke_state : std_logic_vector(1 downto 0);
  signal bombcooke_bombxsample : std_logic_vector(3 downto 0);
  signal bombcooke_bombysample : std_logic_vector(3 downto 0);
  signal bombcookf_state : std_logic_vector(1 downto 0);
  signal bombcookf_bombxsample : std_logic_vector(3 downto 0);
  signal bombcookf_bombysample : std_logic_vector(3 downto 0);
  signal bombcookg_state : std_logic_vector(1 downto 0);
  signal bombcookg_bombxsample : std_logic_vector(3 downto 0);
  signal bombcookg_bombysample : std_logic_vector(3 downto 0);
  signal bombcookh_state : std_logic_vector(1 downto 0);
  signal bombcookh_bombxsample : std_logic_vector(3 downto 0);
  signal bombcookh_bombysample : std_logic_vector(3 downto 0);
  signal mapmech_t28_state : std_logic_vector(1 downto 0);
  signal mapmech_t30_state : std_logic_vector(1 downto 0);
  signal mapmech_t36_state : std_logic_vector(1 downto 0);
  signal mapmech_t37_state : std_logic_vector(1 downto 0);
  signal mapmech_t38_state : std_logic_vector(1 downto 0);
  signal mapmech_t39_state : std_logic_vector(1 downto 0);
  signal mapmech_t40_state : std_logic_vector(1 downto 0);
  signal mapmech_t41_state : std_logic_vector(1 downto 0);
  signal mapmech_t42_state : std_logic_vector(1 downto 0);
  signal mapmech_t46_state : std_logic_vector(1 downto 0);
  signal mapmech_t48_state : std_logic_vector(1 downto 0);
  signal mapmech_t52_state : std_logic_vector(1 downto 0);
  signal mapmech_t54_state : std_logic_vector(1 downto 0);
  signal mapmech_t57_state : std_logic_vector(1 downto 0);
  signal mapmech_t58_state : std_logic_vector(1 downto 0);
  signal mapmech_t59_state : std_logic_vector(1 downto 0);
  signal mapmech_t63_state : std_logic_vector(1 downto 0);
  signal mapmech_t64_state : std_logic_vector(1 downto 0);
  signal mapmech_t65_state : std_logic_vector(1 downto 0);
  signal mapmech_t104_state : std_logic_vector(1 downto 0);
  signal mapmech_t105_state : std_logic_vector(1 downto 0);
  signal mapmech_t68_state : std_logic_vector(1 downto 0);
  signal mapmech_t106_state : std_logic_vector(1 downto 0);
  signal mapmech_t70_state : std_logic_vector(1 downto 0);
  signal mapmech_t74_state : std_logic_vector(1 downto 0);
  signal mapmech_t76_state : std_logic_vector(1 downto 0);
  signal mapmech_t80_state : std_logic_vector(1 downto 0);
  signal mapmech_t81_state : std_logic_vector(1 downto 0);
  signal mapmech_t82_state : std_logic_vector(1 downto 0);
  signal mapmech_t83_state : std_logic_vector(1 downto 0);
  signal mapmech_t84_state : std_logic_vector(1 downto 0);
  signal mapmech_t85_state : std_logic_vector(1 downto 0);
  signal mapmech_t86_state : std_logic_vector(1 downto 0);
  signal mapmech_t16_state : std_logic_vector(1 downto 0);
  signal mapmech_t17_state : std_logic_vector(1 downto 0);
  signal mapmech_t18_state : std_logic_vector(1 downto 0);
  signal mapmech_t92_state : std_logic_vector(1 downto 0);
  signal mapmech_t94_state : std_logic_vector(1 downto 0);
  signal mapmech_t96_state : std_logic_vector(1 downto 0);
  signal mapmech_t26_state : std_logic_vector(1 downto 0);
  signal bombcooka_n_0, bombcooka_n_1, bombcooka_n_2, bombcooka_n_3, bombcooka_n_4 : std_logic;
  signal bombcooka_n_14, bombcookb_n_0, bombcookb_n_1, bombcookb_n_2, bombcookb_n_3 : std_logic;
  signal bombcookb_n_4, bombcookb_n_14, bombcookc_n_0, bombcookc_n_1, bombcookc_n_2 : std_logic;
  signal bombcookc_n_3, bombcookc_n_4, bombcookc_n_14, bombcookd_n_0, bombcookd_n_1 : std_logic;
  signal bombcookd_n_2, bombcookd_n_3, bombcookd_n_4, bombcookd_n_14, bombcooke_n_0 : std_logic;
  signal bombcooke_n_1, bombcooke_n_2, bombcooke_n_3, bombcooke_n_4, bombcooke_n_14 : std_logic;
  signal bombcookf_n_0, bombcookf_n_1, bombcookf_n_2, bombcookf_n_3, bombcookf_n_4 : std_logic;
  signal bombcookf_n_14, bombcookg_n_0, bombcookg_n_1, bombcookg_n_2, bombcookg_n_3 : std_logic;
  signal bombcookg_n_4, bombcookg_n_14, bombcookh_n_0, bombcookh_n_1, bombcookh_n_2 : std_logic;
  signal bombcookh_n_3, bombcookh_n_4, bombcookh_n_14, bombselp1_n_0, bombselp1_n_1 : std_logic;
  signal bombselp1_n_2, bombselp1_n_3, bombselp1_n_4, bombselp1_n_5, bombselp1_n_6 : std_logic;
  signal bombselp1_n_7, bombselp1_n_8, bombselp1_n_12, bombselp2_n_0, bombselp2_n_1 : std_logic;
  signal bombselp2_n_2, bombselp2_n_3, bombselp2_n_4, bombselp2_n_5, bombselp2_n_6 : std_logic;
  signal bombselp2_n_7, bombselp2_n_8, bombselp2_n_12, mapmech_t13_n_0, mapmech_t13_n_1 : std_logic;
  signal mapmech_t13_n_2, mapmech_t13_state, mapmech_t14_n_0, mapmech_t14_n_1, mapmech_t14_n_2 : std_logic;
  signal mapmech_t14_state, mapmech_t15_n_0, mapmech_t15_n_1, mapmech_t15_n_2, mapmech_t15_state : std_logic;
  signal mapmech_t16_n_1, mapmech_t16_n_2, mapmech_t16_n_3, mapmech_t16_n_4, mapmech_t16_n_5 : std_logic;
  signal mapmech_t16_n_6, mapmech_t16_n_7, mapmech_t16_n_8, mapmech_t17_n_1, mapmech_t17_n_2 : std_logic;
  signal mapmech_t17_n_3, mapmech_t17_n_4, mapmech_t17_n_5, mapmech_t17_n_6, mapmech_t17_n_7 : std_logic;
  signal mapmech_t17_n_9, mapmech_t18_n_1, mapmech_t18_n_2, mapmech_t18_n_3, mapmech_t18_n_4 : std_logic;
  signal mapmech_t18_n_5, mapmech_t18_n_6, mapmech_t18_n_7, mapmech_t18_n_8, mapmech_t19_n_0 : std_logic;
  signal mapmech_t19_n_1, mapmech_t19_n_2, mapmech_t19_state, mapmech_t20_n_0, mapmech_t20_n_1 : std_logic;
  signal mapmech_t20_n_2, mapmech_t20_state, mapmech_t21_n_0, mapmech_t21_n_1, mapmech_t21_n_2 : std_logic;
  signal mapmech_t21_state, mapmech_t24_n_0, mapmech_t24_n_1, mapmech_t24_n_2, mapmech_t24_state : std_logic;
  signal mapmech_t26_n_1, mapmech_t26_n_2, mapmech_t26_n_3, mapmech_t26_n_4, mapmech_t26_n_5 : std_logic;
  signal mapmech_t26_n_6, mapmech_t26_n_7, mapmech_t26_n_8, mapmech_t28_n_1, mapmech_t28_n_2 : std_logic;
  signal mapmech_t28_n_3, mapmech_t28_n_4, mapmech_t28_n_5, mapmech_t28_n_6, mapmech_t28_n_7 : std_logic;
  signal mapmech_t28_n_9, mapmech_t30_n_1, mapmech_t30_n_2, mapmech_t30_n_3, mapmech_t30_n_4 : std_logic;
  signal mapmech_t30_n_5, mapmech_t30_n_6, mapmech_t30_n_7, mapmech_t30_n_9, mapmech_t32_n_0 : std_logic;
  signal mapmech_t32_n_1, mapmech_t32_n_2, mapmech_t32_state, mapmech_t35_n_0, mapmech_t35_n_1 : std_logic;
  signal mapmech_t35_n_2, mapmech_t35_state, mapmech_t36_n_1, mapmech_t36_n_2, mapmech_t36_n_3 : std_logic;
  signal mapmech_t36_n_4, mapmech_t36_n_5, mapmech_t36_n_6, mapmech_t36_n_7, mapmech_t36_n_9 : std_logic;
  signal mapmech_t37_n_1, mapmech_t37_n_2, mapmech_t37_n_3, mapmech_t37_n_4, mapmech_t37_n_5 : std_logic;
  signal mapmech_t37_n_6, mapmech_t37_n_7, mapmech_t37_n_8, mapmech_t38_n_1, mapmech_t38_n_2 : std_logic;
  signal mapmech_t38_n_3, mapmech_t38_n_4, mapmech_t38_n_5, mapmech_t38_n_6, mapmech_t38_n_7 : std_logic;
  signal mapmech_t38_n_8, mapmech_t39_n_1, mapmech_t39_n_2, mapmech_t39_n_3, mapmech_t39_n_4 : std_logic;
  signal mapmech_t39_n_5, mapmech_t39_n_6, mapmech_t39_n_7, mapmech_t39_n_9, mapmech_t40_n_1 : std_logic;
  signal mapmech_t40_n_2, mapmech_t40_n_3, mapmech_t40_n_4, mapmech_t40_n_5, mapmech_t40_n_6 : std_logic;
  signal mapmech_t40_n_7, mapmech_t40_n_8, mapmech_t41_n_1, mapmech_t41_n_2, mapmech_t41_n_3 : std_logic;
  signal mapmech_t41_n_4, mapmech_t41_n_5, mapmech_t41_n_6, mapmech_t41_n_7, mapmech_t41_n_8 : std_logic;
  signal mapmech_t42_n_1, mapmech_t42_n_2, mapmech_t42_n_3, mapmech_t42_n_4, mapmech_t42_n_5 : std_logic;
  signal mapmech_t42_n_6, mapmech_t42_n_7, mapmech_t42_n_8, mapmech_t43_n_0, mapmech_t43_n_1 : std_logic;
  signal mapmech_t43_n_2, mapmech_t43_state, mapmech_t46_n_1, mapmech_t46_n_2, mapmech_t46_n_3 : std_logic;
  signal mapmech_t46_n_4, mapmech_t46_n_5, mapmech_t46_n_6, mapmech_t46_n_7, mapmech_t46_n_9 : std_logic;
  signal mapmech_t48_n_1, mapmech_t48_n_2, mapmech_t48_n_3, mapmech_t48_n_4, mapmech_t48_n_5 : std_logic;
  signal mapmech_t48_n_6, mapmech_t48_n_7, mapmech_t48_n_9, mapmech_t50_n_0, mapmech_t50_n_1 : std_logic;
  signal mapmech_t50_n_2, mapmech_t50_state, mapmech_t52_n_1, mapmech_t52_n_2, mapmech_t52_n_3 : std_logic;
  signal mapmech_t52_n_4, mapmech_t52_n_5, mapmech_t52_n_6, mapmech_t52_n_7, mapmech_t52_n_9 : std_logic;
  signal mapmech_t54_n_1, mapmech_t54_n_2, mapmech_t54_n_3, mapmech_t54_n_4, mapmech_t54_n_5 : std_logic;
  signal mapmech_t54_n_6, mapmech_t54_n_7, mapmech_t54_n_8, mapmech_t57_n_1, mapmech_t57_n_2 : std_logic;
  signal mapmech_t57_n_3, mapmech_t57_n_4, mapmech_t57_n_5, mapmech_t57_n_6, mapmech_t57_n_7 : std_logic;
  signal mapmech_t57_n_9, mapmech_t58_n_1, mapmech_t58_n_2, mapmech_t58_n_3, mapmech_t58_n_4 : std_logic;
  signal mapmech_t58_n_5, mapmech_t58_n_6, mapmech_t58_n_7, mapmech_t58_n_8, mapmech_t59_n_1 : std_logic;
  signal mapmech_t59_n_2, mapmech_t59_n_3, mapmech_t59_n_4, mapmech_t59_n_5, mapmech_t59_n_6 : std_logic;
  signal mapmech_t59_n_7, mapmech_t59_n_8, mapmech_t60_n_0, mapmech_t60_n_1, mapmech_t60_n_2 : std_logic;
  signal mapmech_t60_state, mapmech_t61_n_0, mapmech_t61_n_1, mapmech_t61_n_2, mapmech_t61_state : std_logic;
  signal mapmech_t62_n_0, mapmech_t62_n_1, mapmech_t62_n_2, mapmech_t62_state, mapmech_t63_n_1 : std_logic;
  signal mapmech_t63_n_2, mapmech_t63_n_3, mapmech_t63_n_4, mapmech_t63_n_5, mapmech_t63_n_6 : std_logic;
  signal mapmech_t63_n_7, mapmech_t63_n_9, mapmech_t64_n_1, mapmech_t64_n_2, mapmech_t64_n_3 : std_logic;
  signal mapmech_t64_n_4, mapmech_t64_n_5, mapmech_t64_n_6, mapmech_t64_n_7, mapmech_t64_n_9 : std_logic;
  signal mapmech_t65_n_1, mapmech_t65_n_2, mapmech_t65_n_3, mapmech_t65_n_4, mapmech_t65_n_5 : std_logic;
  signal mapmech_t65_n_6, mapmech_t65_n_7, mapmech_t65_n_9, mapmech_t68_n_1, mapmech_t68_n_2 : std_logic;
  signal mapmech_t68_n_3, mapmech_t68_n_4, mapmech_t68_n_5, mapmech_t68_n_6, mapmech_t68_n_7 : std_logic;
  signal mapmech_t68_n_8, mapmech_t70_n_1, mapmech_t70_n_2, mapmech_t70_n_3, mapmech_t70_n_4 : std_logic;
  signal mapmech_t70_n_5, mapmech_t70_n_6, mapmech_t70_n_7, mapmech_t70_n_9, mapmech_t72_n_0 : std_logic;
  signal mapmech_t72_n_1, mapmech_t72_n_2, mapmech_t72_state, mapmech_t74_n_1, mapmech_t74_n_2 : std_logic;
  signal mapmech_t74_n_3, mapmech_t74_n_4, mapmech_t74_n_5, mapmech_t74_n_6, mapmech_t74_n_7 : std_logic;
  signal mapmech_t74_n_9, mapmech_t76_n_1, mapmech_t76_n_2, mapmech_t76_n_3, mapmech_t76_n_4 : std_logic;
  signal mapmech_t76_n_5, mapmech_t76_n_6, mapmech_t76_n_7, mapmech_t76_n_9, mapmech_t79_n_0 : std_logic;
  signal mapmech_t79_n_1, mapmech_t79_n_2, mapmech_t79_state, mapmech_t80_n_1, mapmech_t80_n_2 : std_logic;
  signal mapmech_t80_n_3, mapmech_t80_n_4, mapmech_t80_n_5, mapmech_t80_n_6, mapmech_t80_n_7 : std_logic;
  signal mapmech_t80_n_9, mapmech_t81_n_1, mapmech_t81_n_2, mapmech_t81_n_3, mapmech_t81_n_4 : std_logic;
  signal mapmech_t81_n_5, mapmech_t81_n_6, mapmech_t81_n_7, mapmech_t81_n_8, mapmech_t82_n_1 : std_logic;
  signal mapmech_t82_n_2, mapmech_t82_n_3, mapmech_t82_n_4, mapmech_t82_n_5, mapmech_t82_n_6 : std_logic;
  signal mapmech_t82_n_7, mapmech_t82_n_8, mapmech_t83_n_1, mapmech_t83_n_2, mapmech_t83_n_3 : std_logic;
  signal mapmech_t83_n_4, mapmech_t83_n_5, mapmech_t83_n_6, mapmech_t83_n_7, mapmech_t83_n_8 : std_logic;
  signal mapmech_t84_n_1, mapmech_t84_n_2, mapmech_t84_n_3, mapmech_t84_n_4, mapmech_t84_n_5 : std_logic;
  signal mapmech_t84_n_6, mapmech_t84_n_7, mapmech_t84_n_9, mapmech_t85_n_1, mapmech_t85_n_2 : std_logic;
  signal mapmech_t85_n_3, mapmech_t85_n_4, mapmech_t85_n_5, mapmech_t85_n_6, mapmech_t85_n_7 : std_logic;
  signal mapmech_t85_n_9, mapmech_t86_n_1, mapmech_t86_n_2, mapmech_t86_n_3, mapmech_t86_n_4 : std_logic;
  signal mapmech_t86_n_5, mapmech_t86_n_6, mapmech_t86_n_7, mapmech_t86_n_8, mapmech_t87_n_0 : std_logic;
  signal mapmech_t87_n_1, mapmech_t87_n_2, mapmech_t87_state, mapmech_t90_n_0, mapmech_t90_n_1 : std_logic;
  signal mapmech_t90_n_2, mapmech_t90_state, mapmech_t92_n_1, mapmech_t92_n_2, mapmech_t92_n_3 : std_logic;
  signal mapmech_t92_n_4, mapmech_t92_n_5, mapmech_t92_n_6, mapmech_t92_n_7, mapmech_t92_n_8 : std_logic;
  signal mapmech_t94_n_1, mapmech_t94_n_2, mapmech_t94_n_3, mapmech_t94_n_4, mapmech_t94_n_5 : std_logic;
  signal mapmech_t94_n_6, mapmech_t94_n_7, mapmech_t94_n_8, mapmech_t96_n_1, mapmech_t96_n_2 : std_logic;
  signal mapmech_t96_n_3, mapmech_t96_n_4, mapmech_t96_n_5, mapmech_t96_n_6, mapmech_t96_n_7 : std_logic;
  signal mapmech_t96_n_9, mapmech_t98_n_0, mapmech_t98_n_1, mapmech_t98_n_2, mapmech_t98_state : std_logic;
  signal mapmech_t101_n_0, mapmech_t101_n_1, mapmech_t101_n_2, mapmech_t101_state, mapmech_t102_n_0 : std_logic;
  signal mapmech_t102_n_1, mapmech_t102_n_2, mapmech_t102_state, mapmech_t103_n_0, mapmech_t103_n_1 : std_logic;
  signal mapmech_t103_n_2, mapmech_t103_state, mapmech_t104_n_1, mapmech_t104_n_2, mapmech_t104_n_3 : std_logic;
  signal mapmech_t104_n_4, mapmech_t104_n_5, mapmech_t104_n_6, mapmech_t104_n_7, mapmech_t104_n_9 : std_logic;
  signal mapmech_t105_n_1, mapmech_t105_n_2, mapmech_t105_n_3, mapmech_t105_n_4, mapmech_t105_n_5 : std_logic;
  signal mapmech_t105_n_6, mapmech_t105_n_7, mapmech_t105_n_9, mapmech_t106_n_1, mapmech_t106_n_2 : std_logic;
  signal mapmech_t106_n_3, mapmech_t106_n_4, mapmech_t106_n_5, mapmech_t106_n_6, mapmech_t106_n_7 : std_logic;
  signal mapmech_t106_n_8, mapmech_t107_n_0, mapmech_t107_n_1, mapmech_t107_n_2, mapmech_t107_state : std_logic;
  signal mapmech_t108_n_0, mapmech_t108_n_1, mapmech_t108_n_2, mapmech_t108_state, mapmech_t109_n_0 : std_logic;
  signal mapmech_t109_n_1, mapmech_t109_n_2, mapmech_t109_state, mapmech_xo1, mapmech_xo2 : std_logic;
  signal mapmech_xo3, mapmech_xo4, mapmech_xo5, mapmech_xo6, mapmech_xo7 : std_logic;
  signal mapmech_xo8, mapmech_xo9, mapmech_xyconv_n_1, mapmech_xyconv_n_2, mapmech_xyconv_n_3 : std_logic;
  signal mapmech_xyconv_n_4, mapmech_xyconv_n_5, mapmech_xyconv_n_6, mapmech_xyconv_n_7, mapmech_xyconv_n_8 : std_logic;
  signal mapmech_xyconv_n_10, mapmech_xyconv_n_11, mapmech_xyconv_n_12, mapmech_xyconv_n_14, mapmech_xyconv_n_15 : std_logic;
  signal mapmech_xyconv_n_16, mapmech_yo1, mapmech_yo2, mapmech_yo3, mapmech_yo4 : std_logic;
  signal mapmech_yo5, mapmech_yo6, mapmech_yo7, mapmech_yo8, mapmech_yo9 : std_logic;
  signal n_0, n_105, p1b, p2b : std_logic;

begin

  obstacle_grid(0) <= maptoVGA(241);
  obstacle_grid(1) <= maptoVGA(241);
  obstacle_grid(2) <= maptoVGA(241);
  obstacle_grid(3) <= maptoVGA(241);
  obstacle_grid(4) <= maptoVGA(241);
  obstacle_grid(5) <= maptoVGA(241);
  obstacle_grid(6) <= maptoVGA(241);
  obstacle_grid(7) <= maptoVGA(241);
  obstacle_grid(8) <= maptoVGA(241);
  obstacle_grid(9) <= maptoVGA(241);
  obstacle_grid(10) <= maptoVGA(241);
  obstacle_grid(11) <= maptoVGA(241);
  obstacle_grid(12) <= maptoVGA(217);
  obstacle_grid(13) <= maptoVGA(217);
  obstacle_grid(14) <= maptoVGA(217);
  obstacle_grid(15) <= maptoVGA(31);
  obstacle_grid(16) <= maptoVGA(33);
  obstacle_grid(17) <= maptoVGA(35);
  obstacle_grid(18) <= maptoVGA(217);
  obstacle_grid(19) <= maptoVGA(217);
  obstacle_grid(20) <= maptoVGA(217);
  obstacle_grid(21) <= maptoVGA(241);
  obstacle_grid(22) <= maptoVGA(241);
  obstacle_grid(23) <= maptoVGA(217);
  obstacle_grid(24) <= maptoVGA(241);
  obstacle_grid(25) <= maptoVGA(51);
  obstacle_grid(26) <= maptoVGA(241);
  obstacle_grid(27) <= maptoVGA(55);
  obstacle_grid(28) <= maptoVGA(241);
  obstacle_grid(29) <= maptoVGA(59);
  obstacle_grid(30) <= maptoVGA(241);
  obstacle_grid(31) <= maptoVGA(217);
  obstacle_grid(32) <= maptoVGA(241);
  obstacle_grid(33) <= maptoVGA(241);
  obstacle_grid(34) <= maptoVGA(217);
  obstacle_grid(35) <= maptoVGA(71);
  obstacle_grid(36) <= maptoVGA(73);
  obstacle_grid(37) <= maptoVGA(75);
  obstacle_grid(38) <= maptoVGA(77);
  obstacle_grid(39) <= maptoVGA(79);
  obstacle_grid(40) <= maptoVGA(81);
  obstacle_grid(41) <= maptoVGA(83);
  obstacle_grid(42) <= maptoVGA(217);
  obstacle_grid(43) <= maptoVGA(241);
  obstacle_grid(44) <= maptoVGA(241);
  obstacle_grid(45) <= maptoVGA(91);
  obstacle_grid(46) <= maptoVGA(241);
  obstacle_grid(47) <= maptoVGA(95);
  obstacle_grid(48) <= maptoVGA(241);
  obstacle_grid(49) <= maptoVGA(217);
  obstacle_grid(50) <= maptoVGA(241);
  obstacle_grid(51) <= maptoVGA(103);
  obstacle_grid(52) <= maptoVGA(241);
  obstacle_grid(53) <= maptoVGA(107);
  obstacle_grid(54) <= maptoVGA(241);
  obstacle_grid(55) <= maptoVGA(241);
  obstacle_grid(56) <= maptoVGA(113);
  obstacle_grid(57) <= maptoVGA(115);
  obstacle_grid(58) <= maptoVGA(117);
  obstacle_grid(59) <= maptoVGA(217);
  obstacle_grid(60) <= maptoVGA(217);
  obstacle_grid(61) <= maptoVGA(217);
  obstacle_grid(62) <= maptoVGA(125);
  obstacle_grid(63) <= maptoVGA(127);
  obstacle_grid(64) <= maptoVGA(129);
  obstacle_grid(65) <= maptoVGA(241);
  obstacle_grid(66) <= maptoVGA(241);
  obstacle_grid(67) <= maptoVGA(135);
  obstacle_grid(68) <= maptoVGA(241);
  obstacle_grid(69) <= maptoVGA(139);
  obstacle_grid(70) <= maptoVGA(241);
  obstacle_grid(71) <= maptoVGA(217);
  obstacle_grid(72) <= maptoVGA(241);
  obstacle_grid(73) <= maptoVGA(147);
  obstacle_grid(74) <= maptoVGA(241);
  obstacle_grid(75) <= maptoVGA(151);
  obstacle_grid(76) <= maptoVGA(241);
  obstacle_grid(77) <= maptoVGA(241);
  obstacle_grid(78) <= maptoVGA(217);
  obstacle_grid(79) <= maptoVGA(159);
  obstacle_grid(80) <= maptoVGA(161);
  obstacle_grid(81) <= maptoVGA(163);
  obstacle_grid(82) <= maptoVGA(165);
  obstacle_grid(83) <= maptoVGA(167);
  obstacle_grid(84) <= maptoVGA(169);
  obstacle_grid(85) <= maptoVGA(171);
  obstacle_grid(86) <= maptoVGA(217);
  obstacle_grid(87) <= maptoVGA(241);
  obstacle_grid(88) <= maptoVGA(241);
  obstacle_grid(89) <= maptoVGA(217);
  obstacle_grid(90) <= maptoVGA(241);
  obstacle_grid(91) <= maptoVGA(183);
  obstacle_grid(92) <= maptoVGA(241);
  obstacle_grid(93) <= maptoVGA(187);
  obstacle_grid(94) <= maptoVGA(241);
  obstacle_grid(95) <= maptoVGA(191);
  obstacle_grid(96) <= maptoVGA(241);
  obstacle_grid(97) <= maptoVGA(217);
  obstacle_grid(98) <= maptoVGA(241);
  obstacle_grid(99) <= maptoVGA(241);
  obstacle_grid(100) <= maptoVGA(217);
  obstacle_grid(101) <= maptoVGA(217);
  obstacle_grid(102) <= maptoVGA(217);
  obstacle_grid(103) <= maptoVGA(207);
  obstacle_grid(104) <= maptoVGA(209);
  obstacle_grid(105) <= maptoVGA(211);
  obstacle_grid(106) <= maptoVGA(217);
  obstacle_grid(107) <= maptoVGA(217);
  obstacle_grid(108) <= maptoVGA(217);
  obstacle_grid(109) <= maptoVGA(241);
  obstacle_grid(110) <= maptoVGA(241);
  obstacle_grid(111) <= maptoVGA(241);
  obstacle_grid(112) <= maptoVGA(241);
  obstacle_grid(113) <= maptoVGA(241);
  obstacle_grid(114) <= maptoVGA(241);
  obstacle_grid(115) <= maptoVGA(241);
  obstacle_grid(116) <= maptoVGA(241);
  obstacle_grid(117) <= maptoVGA(241);
  obstacle_grid(118) <= maptoVGA(241);
  obstacle_grid(119) <= maptoVGA(241);
  obstacle_grid(120) <= maptoVGA(241);
  maptoVGA(0) <= maptoVGA(241);
  maptoVGA(1) <= maptoVGA(241);
  maptoVGA(2) <= maptoVGA(241);
  maptoVGA(3) <= maptoVGA(241);
  maptoVGA(4) <= maptoVGA(241);
  maptoVGA(5) <= maptoVGA(241);
  maptoVGA(6) <= maptoVGA(241);
  maptoVGA(7) <= maptoVGA(241);
  maptoVGA(8) <= maptoVGA(241);
  maptoVGA(9) <= maptoVGA(241);
  maptoVGA(10) <= maptoVGA(241);
  maptoVGA(11) <= maptoVGA(241);
  maptoVGA(12) <= maptoVGA(241);
  maptoVGA(13) <= maptoVGA(241);
  maptoVGA(14) <= maptoVGA(241);
  maptoVGA(15) <= maptoVGA(241);
  maptoVGA(16) <= maptoVGA(241);
  maptoVGA(17) <= maptoVGA(241);
  maptoVGA(18) <= maptoVGA(241);
  maptoVGA(19) <= maptoVGA(241);
  maptoVGA(20) <= maptoVGA(241);
  maptoVGA(21) <= maptoVGA(241);
  maptoVGA(22) <= maptoVGA(241);
  maptoVGA(23) <= maptoVGA(241);
  maptoVGA(25) <= maptoVGA(217);
  maptoVGA(27) <= maptoVGA(217);
  maptoVGA(29) <= maptoVGA(217);
  maptoVGA(37) <= maptoVGA(217);
  maptoVGA(39) <= maptoVGA(217);
  maptoVGA(41) <= maptoVGA(217);
  maptoVGA(42) <= maptoVGA(241);
  maptoVGA(43) <= maptoVGA(241);
  maptoVGA(44) <= maptoVGA(241);
  maptoVGA(45) <= maptoVGA(241);
  maptoVGA(47) <= maptoVGA(217);
  maptoVGA(48) <= maptoVGA(241);
  maptoVGA(49) <= maptoVGA(241);
  maptoVGA(52) <= maptoVGA(241);
  maptoVGA(53) <= maptoVGA(241);
  maptoVGA(56) <= maptoVGA(241);
  maptoVGA(57) <= maptoVGA(241);
  maptoVGA(60) <= maptoVGA(241);
  maptoVGA(61) <= maptoVGA(241);
  maptoVGA(63) <= maptoVGA(217);
  maptoVGA(64) <= maptoVGA(241);
  maptoVGA(65) <= maptoVGA(241);
  maptoVGA(66) <= maptoVGA(241);
  maptoVGA(67) <= maptoVGA(241);
  maptoVGA(69) <= maptoVGA(217);
  maptoVGA(85) <= maptoVGA(217);
  maptoVGA(86) <= maptoVGA(241);
  maptoVGA(87) <= maptoVGA(241);
  maptoVGA(88) <= maptoVGA(241);
  maptoVGA(89) <= maptoVGA(241);
  maptoVGA(92) <= maptoVGA(241);
  maptoVGA(93) <= maptoVGA(241);
  maptoVGA(96) <= maptoVGA(241);
  maptoVGA(97) <= maptoVGA(241);
  maptoVGA(99) <= maptoVGA(217);
  maptoVGA(100) <= maptoVGA(241);
  maptoVGA(101) <= maptoVGA(241);
  maptoVGA(104) <= maptoVGA(241);
  maptoVGA(105) <= maptoVGA(241);
  maptoVGA(108) <= maptoVGA(241);
  maptoVGA(109) <= maptoVGA(241);
  maptoVGA(110) <= maptoVGA(241);
  maptoVGA(111) <= maptoVGA(241);
  maptoVGA(119) <= maptoVGA(217);
  maptoVGA(121) <= maptoVGA(217);
  maptoVGA(123) <= maptoVGA(217);
  maptoVGA(130) <= maptoVGA(241);
  maptoVGA(131) <= maptoVGA(241);
  maptoVGA(132) <= maptoVGA(241);
  maptoVGA(133) <= maptoVGA(241);
  maptoVGA(136) <= maptoVGA(241);
  maptoVGA(137) <= maptoVGA(241);
  maptoVGA(140) <= maptoVGA(241);
  maptoVGA(141) <= maptoVGA(241);
  maptoVGA(143) <= maptoVGA(217);
  maptoVGA(144) <= maptoVGA(241);
  maptoVGA(145) <= maptoVGA(241);
  maptoVGA(148) <= maptoVGA(241);
  maptoVGA(149) <= maptoVGA(241);
  maptoVGA(152) <= maptoVGA(241);
  maptoVGA(153) <= maptoVGA(241);
  maptoVGA(154) <= maptoVGA(241);
  maptoVGA(155) <= maptoVGA(241);
  maptoVGA(157) <= maptoVGA(217);
  maptoVGA(173) <= maptoVGA(217);
  maptoVGA(174) <= maptoVGA(241);
  maptoVGA(175) <= maptoVGA(241);
  maptoVGA(176) <= maptoVGA(241);
  maptoVGA(177) <= maptoVGA(241);
  maptoVGA(179) <= maptoVGA(217);
  maptoVGA(180) <= maptoVGA(241);
  maptoVGA(181) <= maptoVGA(241);
  maptoVGA(184) <= maptoVGA(241);
  maptoVGA(185) <= maptoVGA(241);
  maptoVGA(188) <= maptoVGA(241);
  maptoVGA(189) <= maptoVGA(241);
  maptoVGA(192) <= maptoVGA(241);
  maptoVGA(193) <= maptoVGA(241);
  maptoVGA(195) <= maptoVGA(217);
  maptoVGA(196) <= maptoVGA(241);
  maptoVGA(197) <= maptoVGA(241);
  maptoVGA(198) <= maptoVGA(241);
  maptoVGA(199) <= maptoVGA(241);
  maptoVGA(201) <= maptoVGA(217);
  maptoVGA(203) <= maptoVGA(217);
  maptoVGA(205) <= maptoVGA(217);
  maptoVGA(213) <= maptoVGA(217);
  maptoVGA(215) <= maptoVGA(217);
  maptoVGA(218) <= maptoVGA(241);
  maptoVGA(219) <= maptoVGA(241);
  maptoVGA(220) <= maptoVGA(241);
  maptoVGA(221) <= maptoVGA(241);
  maptoVGA(222) <= maptoVGA(241);
  maptoVGA(223) <= maptoVGA(241);
  maptoVGA(224) <= maptoVGA(241);
  maptoVGA(225) <= maptoVGA(241);
  maptoVGA(226) <= maptoVGA(241);
  maptoVGA(227) <= maptoVGA(241);
  maptoVGA(228) <= maptoVGA(241);
  maptoVGA(229) <= maptoVGA(241);
  maptoVGA(230) <= maptoVGA(241);
  maptoVGA(231) <= maptoVGA(241);
  maptoVGA(232) <= maptoVGA(241);
  maptoVGA(233) <= maptoVGA(241);
  maptoVGA(234) <= maptoVGA(241);
  maptoVGA(235) <= maptoVGA(241);
  maptoVGA(236) <= maptoVGA(241);
  maptoVGA(237) <= maptoVGA(241);
  maptoVGA(238) <= maptoVGA(241);
  maptoVGA(239) <= maptoVGA(241);
  maptoVGA(240) <= maptoVGA(241);
  g1 : BUFFD1P5BWP7T port map(I => reset, Z => n_0);
  drc_bufs : BUFFD2BWP7T port map(I => lethal_flag, Z => n_105);
  bombselp1_g181 : INVD0BWP7T port map(I => bombselp1_n_12, ZN => bombselp1_n_6);
  bombselp1_g236 : NR2XD0BWP7T port map(A1 => bombselp1_n_5, A2 => bombselp1_n_7, ZN => bombnop1(3));
  bombselp1_g237 : NR2XD0BWP7T port map(A1 => bombselp1_n_5, A2 => bombselp1_state(2), ZN => bombnop1(1));
  bombselp1_g238 : CKAN2D1BWP7T port map(A1 => bombselp1_n_12, A2 => bombselp1_n_7, Z => bombnop1(0));
  bombselp1_g239 : CKAN2D1BWP7T port map(A1 => bombselp1_n_12, A2 => bombselp1_state(2), Z => bombnop1(2));
  bombselp1_g240 : ND2D1BWP7T port map(A1 => bombselp1_state(1), A2 => bombselp1_state(0), ZN => bombselp1_n_5);
  bombselp1_g241 : INR2XD0BWP7T port map(A1 => bombselp1_state(0), B1 => bombselp1_state(1), ZN => bombselp1_n_12);
  bombselp1_state_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => bombselp1_n_8, D => p1b, Q => bombselp1_state(0));
  bombselp1_g244 : INVD1BWP7T port map(I => reset, ZN => bombselp1_n_8);
  bombselp1_g274 : MOAI22D0BWP7T port map(A1 => bombselp1_n_7, A2 => bombselp1_n_1, B1 => bombselp1_n_2, B2 => bombselp1_n_1, ZN => bombselp1_n_4);
  bombselp1_g275 : OAI22D0BWP7T port map(A1 => bombselp1_n_0, A2 => bombselp1_n_1, B1 => bombselp1_n_6, B2 => p1b, ZN => bombselp1_n_3);
  bombselp1_g276 : MOAI22D0BWP7T port map(A1 => bombselp1_n_0, A2 => bombselp1_state(2), B1 => bombselp1_n_0, B2 => bombselp1_state(2), ZN => bombselp1_n_2);
  bombselp1_g277 : INR2D1BWP7T port map(A1 => bombselp1_state(0), B1 => p1b, ZN => bombselp1_n_1);
  bombselp1_state_reg_2 : DFKCND1BWP7T port map(CP => clk, CN => bombselp1_n_8, D => bombselp1_n_4, Q => bombselp1_state(2), QN => bombselp1_n_7);
  bombselp1_state_reg_1 : DFKCND1BWP7T port map(CP => clk, CN => bombselp1_n_8, D => bombselp1_n_3, Q => bombselp1_state(1), QN => bombselp1_n_0);
  bombselp2_g181 : INVD0BWP7T port map(I => bombselp2_n_12, ZN => bombselp2_n_6);
  bombselp2_g236 : NR2XD0BWP7T port map(A1 => bombselp2_n_5, A2 => bombselp2_n_7, ZN => bombnop2(3));
  bombselp2_g237 : NR2XD0BWP7T port map(A1 => bombselp2_n_5, A2 => bombselp2_state(2), ZN => bombnop2(1));
  bombselp2_g238 : CKAN2D1BWP7T port map(A1 => bombselp2_n_12, A2 => bombselp2_n_7, Z => bombnop2(0));
  bombselp2_g239 : CKAN2D1BWP7T port map(A1 => bombselp2_n_12, A2 => bombselp2_state(2), Z => bombnop2(2));
  bombselp2_g240 : ND2D1BWP7T port map(A1 => bombselp2_state(1), A2 => bombselp2_state(0), ZN => bombselp2_n_5);
  bombselp2_g241 : INR2XD0BWP7T port map(A1 => bombselp2_state(0), B1 => bombselp2_state(1), ZN => bombselp2_n_12);
  bombselp2_state_reg_0 : DFKCNQD1BWP7T port map(CP => clk, CN => bombselp2_n_8, D => p2b, Q => bombselp2_state(0));
  bombselp2_g244 : INVD1BWP7T port map(I => reset, ZN => bombselp2_n_8);
  bombselp2_g274 : MOAI22D0BWP7T port map(A1 => bombselp2_n_7, A2 => bombselp2_n_1, B1 => bombselp2_n_2, B2 => bombselp2_n_1, ZN => bombselp2_n_4);
  bombselp2_g275 : OAI22D0BWP7T port map(A1 => bombselp2_n_0, A2 => bombselp2_n_1, B1 => bombselp2_n_6, B2 => p2b, ZN => bombselp2_n_3);
  bombselp2_g276 : MOAI22D0BWP7T port map(A1 => bombselp2_n_0, A2 => bombselp2_state(2), B1 => bombselp2_n_0, B2 => bombselp2_state(2), ZN => bombselp2_n_2);
  bombselp2_g277 : INR2D1BWP7T port map(A1 => bombselp2_state(0), B1 => p2b, ZN => bombselp2_n_1);
  bombselp2_state_reg_2 : DFKCND1BWP7T port map(CP => clk, CN => bombselp2_n_8, D => bombselp2_n_4, Q => bombselp2_state(2), QN => bombselp2_n_7);
  bombselp2_state_reg_1 : DFKCND1BWP7T port map(CP => clk, CN => bombselp2_n_8, D => bombselp2_n_3, Q => bombselp2_state(1), QN => bombselp2_n_0);
  pbomb_g17 : INR2XD0BWP7T port map(A1 => p_bombplant, B1 => p_bomb, ZN => p1b);
  pbomb_g18 : AN2D1BWP7T port map(A1 => p_bombplant, A2 => p_bomb, Z => p2b);
  bombcooka_g180 : BUFFD4BWP7T port map(I => bombcooka_state(1), Z => bomb_a_cook);
  bombcooka_g234 : AN2D4BWP7T port map(A1 => bombcooka_state(1), A2 => bombcooka_bombxsample(0), Z => bomb_a_x(0));
  bombcooka_g235 : AN2D4BWP7T port map(A1 => bombcooka_state(1), A2 => bombcooka_bombxsample(2), Z => bomb_a_x(2));
  bombcooka_g236 : AN2D4BWP7T port map(A1 => bombcooka_state(1), A2 => bombcooka_bombxsample(3), Z => bomb_a_x(3));
  bombcooka_g237 : AN2D4BWP7T port map(A1 => bombcooka_state(1), A2 => bombcooka_bombysample(0), Z => bomb_a_y(0));
  bombcooka_g238 : AN2D4BWP7T port map(A1 => bombcooka_state(1), A2 => bombcooka_bombysample(2), Z => bomb_a_y(2));
  bombcooka_g239 : AN2D4BWP7T port map(A1 => bombcooka_state(1), A2 => bombcooka_bombxsample(1), Z => bomb_a_x(1));
  bombcooka_g240 : AN2D4BWP7T port map(A1 => bombcooka_state(1), A2 => bombcooka_bombysample(3), Z => bomb_a_y(3));
  bombcooka_g241 : AN2D4BWP7T port map(A1 => bombcooka_state(1), A2 => bombcooka_bombysample(1), Z => bomb_a_y(1));
  bombcooka_bombxsample_reg_2 : LHQD1BWP7T port map(E => bombcooka_n_14, D => p1_x(2), Q => bombcooka_bombxsample(2));
  bombcooka_bombxsample_reg_0 : LHQD1BWP7T port map(E => bombcooka_n_14, D => p1_x(0), Q => bombcooka_bombxsample(0));
  bombcooka_bombysample_reg_0 : LHQD1BWP7T port map(E => bombcooka_n_14, D => p1_y(0), Q => bombcooka_bombysample(0));
  bombcooka_bombysample_reg_3 : LHQD1BWP7T port map(E => bombcooka_n_14, D => p1_y(3), Q => bombcooka_bombysample(3));
  bombcooka_bombxsample_reg_1 : LHQD1BWP7T port map(E => bombcooka_n_14, D => p1_x(1), Q => bombcooka_bombxsample(1));
  bombcooka_bombysample_reg_2 : LHQD1BWP7T port map(E => bombcooka_n_14, D => p1_y(2), Q => bombcooka_bombysample(2));
  bombcooka_bombxsample_reg_3 : LHQD1BWP7T port map(E => bombcooka_n_14, D => p1_x(3), Q => bombcooka_bombxsample(3));
  bombcooka_bombysample_reg_1 : LHQD1BWP7T port map(E => bombcooka_n_14, D => p1_y(1), Q => bombcooka_bombysample(1));
  bombcooka_g250 : INR2D1BWP7T port map(A1 => bombcooka_state(0), B1 => bombcooka_state(1), ZN => bombcooka_n_14);
  bombcooka_state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => bombcooka_n_0, D => bombcooka_n_3, Q => bombcooka_state(1));
  bombcooka_g251 : MOAI22D0BWP7T port map(A1 => bombcooka_n_2, A2 => bombcooka_state(0), B1 => bombcooka_state(1), B2 => expl, ZN => bombcooka_n_4);
  bombcooka_g252 : AO221D0BWP7T port map(A1 => bombcooka_state(0), A2 => expl, B1 => bombcooka_n_1, B2 => bombcooka_state(1), C => bombcooka_n_14, Z => bombcooka_n_3);
  bombcooka_g253 : IND2D1BWP7T port map(A1 => bombcooka_state(1), B1 => bombnop1(0), ZN => bombcooka_n_2);
  bombcooka_g255 : INVD0BWP7T port map(I => reset, ZN => bombcooka_n_0);
  bombcooka_state_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => bombcooka_n_0, D => bombcooka_n_4, Q => bombcooka_state(0), QN => bombcooka_n_1);
  bombcookb_g180 : BUFFD4BWP7T port map(I => bombcookb_state(1), Z => bomb_b_cook);
  bombcookb_g234 : AN2D4BWP7T port map(A1 => bombcookb_state(1), A2 => bombcookb_bombxsample(0), Z => bomb_b_x(0));
  bombcookb_g235 : AN2D4BWP7T port map(A1 => bombcookb_state(1), A2 => bombcookb_bombxsample(2), Z => bomb_b_x(2));
  bombcookb_g236 : AN2D4BWP7T port map(A1 => bombcookb_state(1), A2 => bombcookb_bombxsample(3), Z => bomb_b_x(3));
  bombcookb_g237 : AN2D4BWP7T port map(A1 => bombcookb_state(1), A2 => bombcookb_bombysample(0), Z => bomb_b_y(0));
  bombcookb_g238 : AN2D4BWP7T port map(A1 => bombcookb_state(1), A2 => bombcookb_bombysample(2), Z => bomb_b_y(2));
  bombcookb_g239 : AN2D4BWP7T port map(A1 => bombcookb_state(1), A2 => bombcookb_bombxsample(1), Z => bomb_b_x(1));
  bombcookb_g240 : AN2D4BWP7T port map(A1 => bombcookb_state(1), A2 => bombcookb_bombysample(3), Z => bomb_b_y(3));
  bombcookb_g241 : AN2D4BWP7T port map(A1 => bombcookb_state(1), A2 => bombcookb_bombysample(1), Z => bomb_b_y(1));
  bombcookb_bombxsample_reg_2 : LHQD1BWP7T port map(E => bombcookb_n_14, D => p1_x(2), Q => bombcookb_bombxsample(2));
  bombcookb_bombxsample_reg_0 : LHQD1BWP7T port map(E => bombcookb_n_14, D => p1_x(0), Q => bombcookb_bombxsample(0));
  bombcookb_bombysample_reg_0 : LHQD1BWP7T port map(E => bombcookb_n_14, D => p1_y(0), Q => bombcookb_bombysample(0));
  bombcookb_bombysample_reg_3 : LHQD1BWP7T port map(E => bombcookb_n_14, D => p1_y(3), Q => bombcookb_bombysample(3));
  bombcookb_bombxsample_reg_1 : LHQD1BWP7T port map(E => bombcookb_n_14, D => p1_x(1), Q => bombcookb_bombxsample(1));
  bombcookb_bombysample_reg_2 : LHQD1BWP7T port map(E => bombcookb_n_14, D => p1_y(2), Q => bombcookb_bombysample(2));
  bombcookb_bombxsample_reg_3 : LHQD1BWP7T port map(E => bombcookb_n_14, D => p1_x(3), Q => bombcookb_bombxsample(3));
  bombcookb_bombysample_reg_1 : LHQD1BWP7T port map(E => bombcookb_n_14, D => p1_y(1), Q => bombcookb_bombysample(1));
  bombcookb_g250 : INR2D1BWP7T port map(A1 => bombcookb_state(0), B1 => bombcookb_state(1), ZN => bombcookb_n_14);
  bombcookb_state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => bombcookb_n_0, D => bombcookb_n_3, Q => bombcookb_state(1));
  bombcookb_g251 : MOAI22D0BWP7T port map(A1 => bombcookb_n_2, A2 => bombcookb_state(0), B1 => bombcookb_state(1), B2 => expl, ZN => bombcookb_n_4);
  bombcookb_g252 : AO221D0BWP7T port map(A1 => bombcookb_state(0), A2 => expl, B1 => bombcookb_n_1, B2 => bombcookb_state(1), C => bombcookb_n_14, Z => bombcookb_n_3);
  bombcookb_g253 : IND2D0BWP7T port map(A1 => bombcookb_state(1), B1 => bombnop1(1), ZN => bombcookb_n_2);
  bombcookb_g255 : INVD0BWP7T port map(I => reset, ZN => bombcookb_n_0);
  bombcookb_state_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => bombcookb_n_0, D => bombcookb_n_4, Q => bombcookb_state(0), QN => bombcookb_n_1);
  bombcookc_g180 : BUFFD4BWP7T port map(I => bombcookc_state(1), Z => bomb_c_cook);
  bombcookc_g234 : AN2D4BWP7T port map(A1 => bombcookc_state(1), A2 => bombcookc_bombxsample(0), Z => bomb_c_x(0));
  bombcookc_g235 : AN2D4BWP7T port map(A1 => bombcookc_state(1), A2 => bombcookc_bombxsample(2), Z => bomb_c_x(2));
  bombcookc_g236 : AN2D4BWP7T port map(A1 => bombcookc_state(1), A2 => bombcookc_bombxsample(3), Z => bomb_c_x(3));
  bombcookc_g237 : AN2D4BWP7T port map(A1 => bombcookc_state(1), A2 => bombcookc_bombysample(0), Z => bomb_c_y(0));
  bombcookc_g238 : AN2D4BWP7T port map(A1 => bombcookc_state(1), A2 => bombcookc_bombysample(2), Z => bomb_c_y(2));
  bombcookc_g239 : AN2D4BWP7T port map(A1 => bombcookc_state(1), A2 => bombcookc_bombxsample(1), Z => bomb_c_x(1));
  bombcookc_g240 : AN2D4BWP7T port map(A1 => bombcookc_state(1), A2 => bombcookc_bombysample(3), Z => bomb_c_y(3));
  bombcookc_g241 : AN2D4BWP7T port map(A1 => bombcookc_state(1), A2 => bombcookc_bombysample(1), Z => bomb_c_y(1));
  bombcookc_bombxsample_reg_2 : LHQD1BWP7T port map(E => bombcookc_n_14, D => p1_x(2), Q => bombcookc_bombxsample(2));
  bombcookc_bombxsample_reg_0 : LHQD1BWP7T port map(E => bombcookc_n_14, D => p1_x(0), Q => bombcookc_bombxsample(0));
  bombcookc_bombysample_reg_0 : LHQD1BWP7T port map(E => bombcookc_n_14, D => p1_y(0), Q => bombcookc_bombysample(0));
  bombcookc_bombysample_reg_3 : LHQD1BWP7T port map(E => bombcookc_n_14, D => p1_y(3), Q => bombcookc_bombysample(3));
  bombcookc_bombxsample_reg_1 : LHQD1BWP7T port map(E => bombcookc_n_14, D => p1_x(1), Q => bombcookc_bombxsample(1));
  bombcookc_bombysample_reg_2 : LHQD1BWP7T port map(E => bombcookc_n_14, D => p1_y(2), Q => bombcookc_bombysample(2));
  bombcookc_bombxsample_reg_3 : LHQD1BWP7T port map(E => bombcookc_n_14, D => p1_x(3), Q => bombcookc_bombxsample(3));
  bombcookc_bombysample_reg_1 : LHQD1BWP7T port map(E => bombcookc_n_14, D => p1_y(1), Q => bombcookc_bombysample(1));
  bombcookc_g250 : INR2D1BWP7T port map(A1 => bombcookc_state(0), B1 => bombcookc_state(1), ZN => bombcookc_n_14);
  bombcookc_state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => bombcookc_n_0, D => bombcookc_n_3, Q => bombcookc_state(1));
  bombcookc_g251 : MOAI22D0BWP7T port map(A1 => bombcookc_n_2, A2 => bombcookc_state(0), B1 => bombcookc_state(1), B2 => expl, ZN => bombcookc_n_4);
  bombcookc_g252 : AO221D0BWP7T port map(A1 => bombcookc_state(0), A2 => expl, B1 => bombcookc_n_1, B2 => bombcookc_state(1), C => bombcookc_n_14, Z => bombcookc_n_3);
  bombcookc_g253 : IND2D1BWP7T port map(A1 => bombcookc_state(1), B1 => bombnop1(2), ZN => bombcookc_n_2);
  bombcookc_g255 : INVD0BWP7T port map(I => reset, ZN => bombcookc_n_0);
  bombcookc_state_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => bombcookc_n_0, D => bombcookc_n_4, Q => bombcookc_state(0), QN => bombcookc_n_1);
  bombcookd_g180 : BUFFD4BWP7T port map(I => bombcookd_state(1), Z => bomb_d_cook);
  bombcookd_g234 : AN2D4BWP7T port map(A1 => bombcookd_state(1), A2 => bombcookd_bombxsample(0), Z => bomb_d_x(0));
  bombcookd_g235 : AN2D4BWP7T port map(A1 => bombcookd_state(1), A2 => bombcookd_bombxsample(2), Z => bomb_d_x(2));
  bombcookd_g236 : AN2D4BWP7T port map(A1 => bombcookd_state(1), A2 => bombcookd_bombxsample(3), Z => bomb_d_x(3));
  bombcookd_g237 : AN2D4BWP7T port map(A1 => bombcookd_state(1), A2 => bombcookd_bombysample(0), Z => bomb_d_y(0));
  bombcookd_g238 : AN2D4BWP7T port map(A1 => bombcookd_state(1), A2 => bombcookd_bombysample(2), Z => bomb_d_y(2));
  bombcookd_g239 : AN2D4BWP7T port map(A1 => bombcookd_state(1), A2 => bombcookd_bombxsample(1), Z => bomb_d_x(1));
  bombcookd_g240 : AN2D4BWP7T port map(A1 => bombcookd_state(1), A2 => bombcookd_bombysample(3), Z => bomb_d_y(3));
  bombcookd_g241 : AN2D4BWP7T port map(A1 => bombcookd_state(1), A2 => bombcookd_bombysample(1), Z => bomb_d_y(1));
  bombcookd_bombxsample_reg_2 : LHQD1BWP7T port map(E => bombcookd_n_14, D => p1_x(2), Q => bombcookd_bombxsample(2));
  bombcookd_bombxsample_reg_0 : LHQD1BWP7T port map(E => bombcookd_n_14, D => p1_x(0), Q => bombcookd_bombxsample(0));
  bombcookd_bombysample_reg_0 : LHQD1BWP7T port map(E => bombcookd_n_14, D => p1_y(0), Q => bombcookd_bombysample(0));
  bombcookd_bombysample_reg_3 : LHQD1BWP7T port map(E => bombcookd_n_14, D => p1_y(3), Q => bombcookd_bombysample(3));
  bombcookd_bombxsample_reg_1 : LHQD1BWP7T port map(E => bombcookd_n_14, D => p1_x(1), Q => bombcookd_bombxsample(1));
  bombcookd_bombysample_reg_2 : LHQD1BWP7T port map(E => bombcookd_n_14, D => p1_y(2), Q => bombcookd_bombysample(2));
  bombcookd_bombxsample_reg_3 : LHQD1BWP7T port map(E => bombcookd_n_14, D => p1_x(3), Q => bombcookd_bombxsample(3));
  bombcookd_bombysample_reg_1 : LHQD1BWP7T port map(E => bombcookd_n_14, D => p1_y(1), Q => bombcookd_bombysample(1));
  bombcookd_g250 : INR2D1BWP7T port map(A1 => bombcookd_state(0), B1 => bombcookd_state(1), ZN => bombcookd_n_14);
  bombcookd_state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => bombcookd_n_0, D => bombcookd_n_3, Q => bombcookd_state(1));
  bombcookd_g251 : MOAI22D0BWP7T port map(A1 => bombcookd_n_2, A2 => bombcookd_state(0), B1 => bombcookd_state(1), B2 => expl, ZN => bombcookd_n_4);
  bombcookd_g252 : AO221D0BWP7T port map(A1 => bombcookd_state(0), A2 => expl, B1 => bombcookd_n_1, B2 => bombcookd_state(1), C => bombcookd_n_14, Z => bombcookd_n_3);
  bombcookd_g253 : IND2D0BWP7T port map(A1 => bombcookd_state(1), B1 => bombnop1(3), ZN => bombcookd_n_2);
  bombcookd_g255 : INVD0BWP7T port map(I => reset, ZN => bombcookd_n_0);
  bombcookd_state_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => bombcookd_n_0, D => bombcookd_n_4, Q => bombcookd_state(0), QN => bombcookd_n_1);
  bombcooke_g180 : BUFFD4BWP7T port map(I => bombcooke_state(1), Z => bomb_e_cook);
  bombcooke_g234 : AN2D4BWP7T port map(A1 => bombcooke_state(1), A2 => bombcooke_bombxsample(0), Z => bomb_e_x(0));
  bombcooke_g235 : AN2D4BWP7T port map(A1 => bombcooke_state(1), A2 => bombcooke_bombxsample(2), Z => bomb_e_x(2));
  bombcooke_g236 : AN2D4BWP7T port map(A1 => bombcooke_state(1), A2 => bombcooke_bombxsample(3), Z => bomb_e_x(3));
  bombcooke_g237 : AN2D4BWP7T port map(A1 => bombcooke_state(1), A2 => bombcooke_bombysample(0), Z => bomb_e_y(0));
  bombcooke_g238 : AN2D4BWP7T port map(A1 => bombcooke_state(1), A2 => bombcooke_bombysample(2), Z => bomb_e_y(2));
  bombcooke_g239 : AN2D4BWP7T port map(A1 => bombcooke_state(1), A2 => bombcooke_bombxsample(1), Z => bomb_e_x(1));
  bombcooke_g240 : AN2D4BWP7T port map(A1 => bombcooke_state(1), A2 => bombcooke_bombysample(3), Z => bomb_e_y(3));
  bombcooke_g241 : AN2D4BWP7T port map(A1 => bombcooke_state(1), A2 => bombcooke_bombysample(1), Z => bomb_e_y(1));
  bombcooke_bombxsample_reg_2 : LHQD1BWP7T port map(E => bombcooke_n_14, D => p2_x(2), Q => bombcooke_bombxsample(2));
  bombcooke_bombxsample_reg_0 : LHQD1BWP7T port map(E => bombcooke_n_14, D => p2_x(0), Q => bombcooke_bombxsample(0));
  bombcooke_bombysample_reg_0 : LHQD1BWP7T port map(E => bombcooke_n_14, D => p2_y(0), Q => bombcooke_bombysample(0));
  bombcooke_bombysample_reg_3 : LHQD1BWP7T port map(E => bombcooke_n_14, D => p2_y(3), Q => bombcooke_bombysample(3));
  bombcooke_bombxsample_reg_1 : LHQD1BWP7T port map(E => bombcooke_n_14, D => p2_x(1), Q => bombcooke_bombxsample(1));
  bombcooke_bombysample_reg_2 : LHQD1BWP7T port map(E => bombcooke_n_14, D => p2_y(2), Q => bombcooke_bombysample(2));
  bombcooke_bombxsample_reg_3 : LHQD1BWP7T port map(E => bombcooke_n_14, D => p2_x(3), Q => bombcooke_bombxsample(3));
  bombcooke_bombysample_reg_1 : LHQD1BWP7T port map(E => bombcooke_n_14, D => p2_y(1), Q => bombcooke_bombysample(1));
  bombcooke_g250 : INR2D1BWP7T port map(A1 => bombcooke_state(0), B1 => bombcooke_state(1), ZN => bombcooke_n_14);
  bombcooke_state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => bombcooke_n_0, D => bombcooke_n_3, Q => bombcooke_state(1));
  bombcooke_g251 : MOAI22D0BWP7T port map(A1 => bombcooke_n_2, A2 => bombcooke_state(0), B1 => bombcooke_state(1), B2 => expl, ZN => bombcooke_n_4);
  bombcooke_g252 : AO221D0BWP7T port map(A1 => bombcooke_state(0), A2 => expl, B1 => bombcooke_n_1, B2 => bombcooke_state(1), C => bombcooke_n_14, Z => bombcooke_n_3);
  bombcooke_g253 : IND2D1BWP7T port map(A1 => bombcooke_state(1), B1 => bombnop2(0), ZN => bombcooke_n_2);
  bombcooke_g255 : INVD0BWP7T port map(I => reset, ZN => bombcooke_n_0);
  bombcooke_state_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => bombcooke_n_0, D => bombcooke_n_4, Q => bombcooke_state(0), QN => bombcooke_n_1);
  bombcookf_g180 : BUFFD4BWP7T port map(I => bombcookf_state(1), Z => bomb_f_cook);
  bombcookf_g234 : AN2D4BWP7T port map(A1 => bombcookf_state(1), A2 => bombcookf_bombxsample(0), Z => bomb_f_x(0));
  bombcookf_g235 : AN2D4BWP7T port map(A1 => bombcookf_state(1), A2 => bombcookf_bombxsample(2), Z => bomb_f_x(2));
  bombcookf_g236 : AN2D4BWP7T port map(A1 => bombcookf_state(1), A2 => bombcookf_bombxsample(3), Z => bomb_f_x(3));
  bombcookf_g237 : AN2D4BWP7T port map(A1 => bombcookf_state(1), A2 => bombcookf_bombysample(0), Z => bomb_f_y(0));
  bombcookf_g238 : AN2D4BWP7T port map(A1 => bombcookf_state(1), A2 => bombcookf_bombysample(2), Z => bomb_f_y(2));
  bombcookf_g239 : AN2D4BWP7T port map(A1 => bombcookf_state(1), A2 => bombcookf_bombxsample(1), Z => bomb_f_x(1));
  bombcookf_g240 : AN2D4BWP7T port map(A1 => bombcookf_state(1), A2 => bombcookf_bombysample(3), Z => bomb_f_y(3));
  bombcookf_g241 : AN2D4BWP7T port map(A1 => bombcookf_state(1), A2 => bombcookf_bombysample(1), Z => bomb_f_y(1));
  bombcookf_bombxsample_reg_2 : LHQD1BWP7T port map(E => bombcookf_n_14, D => p2_x(2), Q => bombcookf_bombxsample(2));
  bombcookf_bombxsample_reg_0 : LHQD1BWP7T port map(E => bombcookf_n_14, D => p2_x(0), Q => bombcookf_bombxsample(0));
  bombcookf_bombysample_reg_0 : LHQD1BWP7T port map(E => bombcookf_n_14, D => p2_y(0), Q => bombcookf_bombysample(0));
  bombcookf_bombysample_reg_3 : LHQD1BWP7T port map(E => bombcookf_n_14, D => p2_y(3), Q => bombcookf_bombysample(3));
  bombcookf_bombxsample_reg_1 : LHQD1BWP7T port map(E => bombcookf_n_14, D => p2_x(1), Q => bombcookf_bombxsample(1));
  bombcookf_bombysample_reg_2 : LHQD1BWP7T port map(E => bombcookf_n_14, D => p2_y(2), Q => bombcookf_bombysample(2));
  bombcookf_bombxsample_reg_3 : LHQD1BWP7T port map(E => bombcookf_n_14, D => p2_x(3), Q => bombcookf_bombxsample(3));
  bombcookf_bombysample_reg_1 : LHQD1BWP7T port map(E => bombcookf_n_14, D => p2_y(1), Q => bombcookf_bombysample(1));
  bombcookf_g250 : INR2D1BWP7T port map(A1 => bombcookf_state(0), B1 => bombcookf_state(1), ZN => bombcookf_n_14);
  bombcookf_state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => bombcookf_n_0, D => bombcookf_n_3, Q => bombcookf_state(1));
  bombcookf_g251 : MOAI22D0BWP7T port map(A1 => bombcookf_n_2, A2 => bombcookf_state(0), B1 => bombcookf_state(1), B2 => expl, ZN => bombcookf_n_4);
  bombcookf_g252 : AO221D0BWP7T port map(A1 => bombcookf_state(0), A2 => expl, B1 => bombcookf_n_1, B2 => bombcookf_state(1), C => bombcookf_n_14, Z => bombcookf_n_3);
  bombcookf_g253 : IND2D0BWP7T port map(A1 => bombcookf_state(1), B1 => bombnop2(1), ZN => bombcookf_n_2);
  bombcookf_g255 : INVD0BWP7T port map(I => reset, ZN => bombcookf_n_0);
  bombcookf_state_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => bombcookf_n_0, D => bombcookf_n_4, Q => bombcookf_state(0), QN => bombcookf_n_1);
  bombcookg_g180 : BUFFD4BWP7T port map(I => bombcookg_state(1), Z => bomb_g_cook);
  bombcookg_g234 : AN2D4BWP7T port map(A1 => bombcookg_state(1), A2 => bombcookg_bombxsample(0), Z => bomb_g_x(0));
  bombcookg_g235 : AN2D4BWP7T port map(A1 => bombcookg_state(1), A2 => bombcookg_bombxsample(2), Z => bomb_g_x(2));
  bombcookg_g236 : AN2D4BWP7T port map(A1 => bombcookg_state(1), A2 => bombcookg_bombxsample(3), Z => bomb_g_x(3));
  bombcookg_g237 : AN2D4BWP7T port map(A1 => bombcookg_state(1), A2 => bombcookg_bombysample(0), Z => bomb_g_y(0));
  bombcookg_g238 : AN2D4BWP7T port map(A1 => bombcookg_state(1), A2 => bombcookg_bombysample(2), Z => bomb_g_y(2));
  bombcookg_g239 : AN2D4BWP7T port map(A1 => bombcookg_state(1), A2 => bombcookg_bombxsample(1), Z => bomb_g_x(1));
  bombcookg_g240 : AN2D4BWP7T port map(A1 => bombcookg_state(1), A2 => bombcookg_bombysample(3), Z => bomb_g_y(3));
  bombcookg_g241 : AN2D4BWP7T port map(A1 => bombcookg_state(1), A2 => bombcookg_bombysample(1), Z => bomb_g_y(1));
  bombcookg_bombxsample_reg_2 : LHQD1BWP7T port map(E => bombcookg_n_14, D => p2_x(2), Q => bombcookg_bombxsample(2));
  bombcookg_bombxsample_reg_0 : LHQD1BWP7T port map(E => bombcookg_n_14, D => p2_x(0), Q => bombcookg_bombxsample(0));
  bombcookg_bombysample_reg_0 : LHQD1BWP7T port map(E => bombcookg_n_14, D => p2_y(0), Q => bombcookg_bombysample(0));
  bombcookg_bombysample_reg_3 : LHQD1BWP7T port map(E => bombcookg_n_14, D => p2_y(3), Q => bombcookg_bombysample(3));
  bombcookg_bombxsample_reg_1 : LHQD1BWP7T port map(E => bombcookg_n_14, D => p2_x(1), Q => bombcookg_bombxsample(1));
  bombcookg_bombysample_reg_2 : LHQD1BWP7T port map(E => bombcookg_n_14, D => p2_y(2), Q => bombcookg_bombysample(2));
  bombcookg_bombxsample_reg_3 : LHQD1BWP7T port map(E => bombcookg_n_14, D => p2_x(3), Q => bombcookg_bombxsample(3));
  bombcookg_bombysample_reg_1 : LHQD1BWP7T port map(E => bombcookg_n_14, D => p2_y(1), Q => bombcookg_bombysample(1));
  bombcookg_g250 : INR2D1BWP7T port map(A1 => bombcookg_state(0), B1 => bombcookg_state(1), ZN => bombcookg_n_14);
  bombcookg_state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => bombcookg_n_0, D => bombcookg_n_3, Q => bombcookg_state(1));
  bombcookg_g251 : MOAI22D0BWP7T port map(A1 => bombcookg_n_2, A2 => bombcookg_state(0), B1 => bombcookg_state(1), B2 => expl, ZN => bombcookg_n_4);
  bombcookg_g252 : AO221D0BWP7T port map(A1 => bombcookg_state(0), A2 => expl, B1 => bombcookg_n_1, B2 => bombcookg_state(1), C => bombcookg_n_14, Z => bombcookg_n_3);
  bombcookg_g253 : IND2D1BWP7T port map(A1 => bombcookg_state(1), B1 => bombnop2(2), ZN => bombcookg_n_2);
  bombcookg_g255 : INVD0BWP7T port map(I => reset, ZN => bombcookg_n_0);
  bombcookg_state_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => bombcookg_n_0, D => bombcookg_n_4, Q => bombcookg_state(0), QN => bombcookg_n_1);
  bombcookh_g180 : BUFFD4BWP7T port map(I => bombcookh_state(1), Z => bomb_h_cook);
  bombcookh_g234 : AN2D4BWP7T port map(A1 => bombcookh_state(1), A2 => bombcookh_bombxsample(0), Z => bomb_h_x(0));
  bombcookh_g235 : AN2D4BWP7T port map(A1 => bombcookh_state(1), A2 => bombcookh_bombxsample(2), Z => bomb_h_x(2));
  bombcookh_g236 : AN2D4BWP7T port map(A1 => bombcookh_state(1), A2 => bombcookh_bombxsample(3), Z => bomb_h_x(3));
  bombcookh_g237 : AN2D4BWP7T port map(A1 => bombcookh_state(1), A2 => bombcookh_bombysample(0), Z => bomb_h_y(0));
  bombcookh_g238 : AN2D4BWP7T port map(A1 => bombcookh_state(1), A2 => bombcookh_bombysample(2), Z => bomb_h_y(2));
  bombcookh_g239 : AN2D4BWP7T port map(A1 => bombcookh_state(1), A2 => bombcookh_bombxsample(1), Z => bomb_h_x(1));
  bombcookh_g240 : AN2D4BWP7T port map(A1 => bombcookh_state(1), A2 => bombcookh_bombysample(3), Z => bomb_h_y(3));
  bombcookh_g241 : AN2D4BWP7T port map(A1 => bombcookh_state(1), A2 => bombcookh_bombysample(1), Z => bomb_h_y(1));
  bombcookh_bombxsample_reg_2 : LHQD1BWP7T port map(E => bombcookh_n_14, D => p2_x(2), Q => bombcookh_bombxsample(2));
  bombcookh_bombxsample_reg_0 : LHQD1BWP7T port map(E => bombcookh_n_14, D => p2_x(0), Q => bombcookh_bombxsample(0));
  bombcookh_bombysample_reg_0 : LHQD1BWP7T port map(E => bombcookh_n_14, D => p2_y(0), Q => bombcookh_bombysample(0));
  bombcookh_bombysample_reg_3 : LHQD1BWP7T port map(E => bombcookh_n_14, D => p2_y(3), Q => bombcookh_bombysample(3));
  bombcookh_bombxsample_reg_1 : LHQD1BWP7T port map(E => bombcookh_n_14, D => p2_x(1), Q => bombcookh_bombxsample(1));
  bombcookh_bombysample_reg_2 : LHQD1BWP7T port map(E => bombcookh_n_14, D => p2_y(2), Q => bombcookh_bombysample(2));
  bombcookh_bombxsample_reg_3 : LHQD1BWP7T port map(E => bombcookh_n_14, D => p2_x(3), Q => bombcookh_bombxsample(3));
  bombcookh_bombysample_reg_1 : LHQD1BWP7T port map(E => bombcookh_n_14, D => p2_y(1), Q => bombcookh_bombysample(1));
  bombcookh_g250 : INR2D1BWP7T port map(A1 => bombcookh_state(0), B1 => bombcookh_state(1), ZN => bombcookh_n_14);
  bombcookh_state_reg_1 : DFKCNQD1BWP7T port map(CP => clk, CN => bombcookh_n_0, D => bombcookh_n_3, Q => bombcookh_state(1));
  bombcookh_g251 : MOAI22D0BWP7T port map(A1 => bombcookh_n_2, A2 => bombcookh_state(0), B1 => bombcookh_state(1), B2 => expl, ZN => bombcookh_n_4);
  bombcookh_g252 : AO221D0BWP7T port map(A1 => bombcookh_state(0), A2 => expl, B1 => bombcookh_n_1, B2 => bombcookh_state(1), C => bombcookh_n_14, Z => bombcookh_n_3);
  bombcookh_g253 : IND2D0BWP7T port map(A1 => bombcookh_state(1), B1 => bombnop2(3), ZN => bombcookh_n_2);
  bombcookh_g255 : INVD0BWP7T port map(I => reset, ZN => bombcookh_n_0);
  bombcookh_state_reg_0 : DFKCND1BWP7T port map(CP => clk, CN => bombcookh_n_0, D => bombcookh_n_4, Q => bombcookh_state(0), QN => bombcookh_n_1);
  mapmech_t98_g68 : INVD4BWP7T port map(I => mapmech_t98_state, ZN => maptoVGA(46));
  mapmech_t98_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t98_n_2, Q => mapmech_t98_state);
  mapmech_t98_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(46), A2 => mapmech_t98_n_1, B => n_0, C => mapmech_t98_n_0, ZN => mapmech_t98_n_2);
  mapmech_t98_g119 : ND2D0BWP7T port map(A1 => mapmech_xo9, A2 => mapmech_yo8, ZN => mapmech_t98_n_1);
  mapmech_t98_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t98_n_0);
  mapmech_t28_g136 : BUFFD4BWP7T port map(I => mapmech_t28_state(1), Z => maptoVGA(186));
  mapmech_t28_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t28_n_7, A2 => mapmech_t28_n_9, Z => maptoVGA(187));
  mapmech_t28_g185 : NR2XD0BWP7T port map(A1 => mapmech_t28_n_4, A2 => n_0, ZN => mapmech_t28_n_6);
  mapmech_t28_g186 : AOI21D0BWP7T port map(A1 => mapmech_t28_n_2, A2 => mapmech_t28_n_3, B => n_0, ZN => mapmech_t28_n_5);
  mapmech_t28_g187 : AOI22D0BWP7T port map(A1 => mapmech_t28_state(1), A2 => mapmech_t28_n_3, B1 => mapmech_t28_state(0), B2 => mapmech_t28_n_1, ZN => mapmech_t28_n_4);
  mapmech_t28_g188 : ND3D0BWP7T port map(A1 => mapmech_xo5, A2 => mapmech_yo2, A3 => n_105, ZN => mapmech_t28_n_3);
  mapmech_t28_g189 : ND2D1BWP7T port map(A1 => mapmech_t28_state(0), A2 => n_105, ZN => mapmech_t28_n_2);
  mapmech_t28_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t28_n_1);
  mapmech_t28_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t28_n_5, Q => mapmech_t28_state(0), QN => mapmech_t28_n_9);
  mapmech_t28_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t28_n_6, Q => mapmech_t28_state(1), QN => mapmech_t28_n_7);
  mapmech_t30_g136 : BUFFD4BWP7T port map(I => mapmech_t30_state(1), Z => maptoVGA(182));
  mapmech_t30_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t30_n_7, A2 => mapmech_t30_n_9, Z => maptoVGA(183));
  mapmech_t30_g185 : NR2XD0BWP7T port map(A1 => mapmech_t30_n_4, A2 => n_0, ZN => mapmech_t30_n_6);
  mapmech_t30_g186 : AOI21D0BWP7T port map(A1 => mapmech_t30_n_2, A2 => mapmech_t30_n_3, B => n_0, ZN => mapmech_t30_n_5);
  mapmech_t30_g187 : AOI22D0BWP7T port map(A1 => mapmech_t30_state(1), A2 => mapmech_t30_n_3, B1 => mapmech_t30_state(0), B2 => mapmech_t30_n_1, ZN => mapmech_t30_n_4);
  mapmech_t30_g188 : ND3D0BWP7T port map(A1 => mapmech_xo7, A2 => mapmech_yo2, A3 => n_105, ZN => mapmech_t30_n_3);
  mapmech_t30_g189 : ND2D1BWP7T port map(A1 => mapmech_t30_state(0), A2 => n_105, ZN => mapmech_t30_n_2);
  mapmech_t30_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t30_n_1);
  mapmech_t30_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t30_n_5, Q => mapmech_t30_state(0), QN => mapmech_t30_n_9);
  mapmech_t30_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t30_n_6, Q => mapmech_t30_state(1), QN => mapmech_t30_n_7);
  mapmech_t32_g68 : INVD4BWP7T port map(I => mapmech_t32_state, ZN => maptoVGA(178));
  mapmech_t32_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t32_n_2, Q => mapmech_t32_state);
  mapmech_t32_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(178), A2 => mapmech_t32_n_1, B => n_0, C => mapmech_t32_n_0, ZN => mapmech_t32_n_2);
  mapmech_t32_g119 : ND2D0BWP7T port map(A1 => mapmech_xo9, A2 => mapmech_yo2, ZN => mapmech_t32_n_1);
  mapmech_t32_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t32_n_0);
  mapmech_t35_g68 : INVD4BWP7T port map(I => mapmech_t35_state, ZN => maptoVGA(172));
  mapmech_t35_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t35_n_2, Q => mapmech_t35_state);
  mapmech_t35_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(172), A2 => mapmech_t35_n_1, B => n_0, C => mapmech_t35_n_0, ZN => mapmech_t35_n_2);
  mapmech_t35_g119 : ND2D0BWP7T port map(A1 => mapmech_yo3, A2 => mapmech_xo1, ZN => mapmech_t35_n_1);
  mapmech_t35_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t35_n_0);
  mapmech_t36_g136 : BUFFD4BWP7T port map(I => mapmech_t36_state(1), Z => maptoVGA(170));
  mapmech_t36_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t36_n_7, A2 => mapmech_t36_n_9, Z => maptoVGA(171));
  mapmech_t36_g185 : NR2XD0BWP7T port map(A1 => mapmech_t36_n_4, A2 => n_0, ZN => mapmech_t36_n_6);
  mapmech_t36_g186 : AOI21D0BWP7T port map(A1 => mapmech_t36_n_2, A2 => mapmech_t36_n_3, B => n_0, ZN => mapmech_t36_n_5);
  mapmech_t36_g187 : AOI22D0BWP7T port map(A1 => mapmech_t36_state(1), A2 => mapmech_t36_n_3, B1 => mapmech_t36_state(0), B2 => mapmech_t36_n_1, ZN => mapmech_t36_n_4);
  mapmech_t36_g188 : ND3D0BWP7T port map(A1 => mapmech_yo3, A2 => mapmech_xo2, A3 => n_105, ZN => mapmech_t36_n_3);
  mapmech_t36_g189 : ND2D1BWP7T port map(A1 => mapmech_t36_state(0), A2 => n_105, ZN => mapmech_t36_n_2);
  mapmech_t36_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t36_n_1);
  mapmech_t36_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t36_n_5, Q => mapmech_t36_state(0), QN => mapmech_t36_n_9);
  mapmech_t36_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t36_n_6, Q => mapmech_t36_state(1), QN => mapmech_t36_n_7);
  mapmech_t37_g135 : BUFFD4BWP7T port map(I => mapmech_t37_state(1), Z => maptoVGA(168));
  mapmech_t37_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t37_n_7, A2 => mapmech_t37_n_8, Z => maptoVGA(169));
  mapmech_t37_g185 : NR2XD0BWP7T port map(A1 => mapmech_t37_n_4, A2 => n_0, ZN => mapmech_t37_n_6);
  mapmech_t37_g186 : AOI21D0BWP7T port map(A1 => mapmech_t37_n_2, A2 => mapmech_t37_n_3, B => n_0, ZN => mapmech_t37_n_5);
  mapmech_t37_g187 : AOI22D0BWP7T port map(A1 => mapmech_t37_state(1), A2 => mapmech_t37_n_3, B1 => mapmech_t37_state(0), B2 => mapmech_t37_n_1, ZN => mapmech_t37_n_4);
  mapmech_t37_g188 : ND3D0BWP7T port map(A1 => mapmech_xo3, A2 => mapmech_yo3, A3 => n_105, ZN => mapmech_t37_n_3);
  mapmech_t37_g189 : ND2D1BWP7T port map(A1 => mapmech_t37_state(0), A2 => n_105, ZN => mapmech_t37_n_2);
  mapmech_t37_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t37_n_1);
  mapmech_t37_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t37_n_5, Q => mapmech_t37_state(0), QN => mapmech_t37_n_8);
  mapmech_t37_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t37_n_6, Q => mapmech_t37_state(1), QN => mapmech_t37_n_7);
  mapmech_xyconv_g491 : INR2XD0BWP7T port map(A1 => lethaltile_x(1), B1 => mapmech_xyconv_n_16, ZN => mapmech_xo7);
  mapmech_xyconv_g492 : NR2XD0BWP7T port map(A1 => mapmech_xyconv_n_16, A2 => lethaltile_x(1), ZN => mapmech_xo5);
  mapmech_xyconv_g493 : INR2XD0BWP7T port map(A1 => lethaltile_x(1), B1 => mapmech_xyconv_n_10, ZN => mapmech_xo6);
  mapmech_xyconv_g494 : NR2XD0BWP7T port map(A1 => mapmech_xyconv_n_11, A2 => lethaltile_y(1), ZN => mapmech_yo4);
  mapmech_xyconv_g495 : NR2XD0BWP7T port map(A1 => mapmech_xyconv_n_10, A2 => lethaltile_x(1), ZN => mapmech_xo4);
  mapmech_xyconv_g496 : NR2XD0BWP7T port map(A1 => mapmech_xyconv_n_12, A2 => lethaltile_y(1), ZN => mapmech_yo5);
  mapmech_xyconv_g497 : INR2XD0BWP7T port map(A1 => lethaltile_y(1), B1 => mapmech_xyconv_n_11, ZN => mapmech_yo6);
  mapmech_xyconv_g498 : NR2XD0BWP7T port map(A1 => mapmech_xyconv_n_15, A2 => lethaltile_x(0), ZN => mapmech_xo8);
  mapmech_xyconv_g499 : NR3D0BWP7T port map(A1 => mapmech_xyconv_n_3, A2 => lethaltile_y(2), A3 => mapmech_xyconv_n_1, ZN => mapmech_yo3);
  mapmech_xyconv_g500 : NR2XD0BWP7T port map(A1 => mapmech_xyconv_n_14, A2 => lethaltile_y(0), ZN => mapmech_yo8);
  mapmech_xyconv_g501 : INR2XD0BWP7T port map(A1 => lethaltile_y(0), B1 => mapmech_xyconv_n_14, ZN => mapmech_yo9);
  mapmech_xyconv_g502 : INR2XD0BWP7T port map(A1 => lethaltile_x(0), B1 => mapmech_xyconv_n_15, ZN => mapmech_xo9);
  mapmech_xyconv_g503 : INR2XD0BWP7T port map(A1 => lethaltile_y(1), B1 => mapmech_xyconv_n_12, ZN => mapmech_yo7);
  mapmech_xyconv_g504 : NR3D0BWP7T port map(A1 => mapmech_xyconv_n_6, A2 => lethaltile_x(2), A3 => mapmech_xyconv_n_2, ZN => mapmech_xo2);
  mapmech_xyconv_g505 : NR3D0BWP7T port map(A1 => mapmech_xyconv_n_4, A2 => lethaltile_x(2), A3 => mapmech_xyconv_n_2, ZN => mapmech_xo3);
  mapmech_xyconv_g506 : NR3D0BWP7T port map(A1 => mapmech_xyconv_n_8, A2 => lethaltile_y(2), A3 => mapmech_xyconv_n_1, ZN => mapmech_yo2);
  mapmech_xyconv_g507 : INR2XD0BWP7T port map(A1 => mapmech_xyconv_n_5, B1 => mapmech_xyconv_n_4, ZN => mapmech_xo1);
  mapmech_xyconv_g508 : IND2D1BWP7T port map(A1 => mapmech_xyconv_n_4, B1 => lethaltile_x(2), ZN => mapmech_xyconv_n_16);
  mapmech_xyconv_g509 : ND2D1BWP7T port map(A1 => mapmech_xyconv_n_5, A2 => lethaltile_x(3), ZN => mapmech_xyconv_n_15);
  mapmech_xyconv_g510 : ND2D1BWP7T port map(A1 => mapmech_xyconv_n_7, A2 => lethaltile_y(3), ZN => mapmech_xyconv_n_14);
  mapmech_xyconv_g511 : INR2XD0BWP7T port map(A1 => mapmech_xyconv_n_7, B1 => mapmech_xyconv_n_3, ZN => mapmech_yo1);
  mapmech_xyconv_g512 : IND2D1BWP7T port map(A1 => mapmech_xyconv_n_3, B1 => lethaltile_y(2), ZN => mapmech_xyconv_n_12);
  mapmech_xyconv_g513 : IND2D1BWP7T port map(A1 => mapmech_xyconv_n_8, B1 => lethaltile_y(2), ZN => mapmech_xyconv_n_11);
  mapmech_xyconv_g514 : IND2D1BWP7T port map(A1 => mapmech_xyconv_n_6, B1 => lethaltile_x(2), ZN => mapmech_xyconv_n_10);
  mapmech_xyconv_g515 : OR2D1BWP7T port map(A1 => lethaltile_y(3), A2 => lethaltile_y(0), Z => mapmech_xyconv_n_8);
  mapmech_xyconv_g516 : NR2XD0BWP7T port map(A1 => lethaltile_y(1), A2 => lethaltile_y(2), ZN => mapmech_xyconv_n_7);
  mapmech_xyconv_g517 : OR2D1BWP7T port map(A1 => lethaltile_x(3), A2 => lethaltile_x(0), Z => mapmech_xyconv_n_6);
  mapmech_xyconv_g518 : NR2XD0BWP7T port map(A1 => lethaltile_x(1), A2 => lethaltile_x(2), ZN => mapmech_xyconv_n_5);
  mapmech_xyconv_g519 : IND2D1BWP7T port map(A1 => lethaltile_x(3), B1 => lethaltile_x(0), ZN => mapmech_xyconv_n_4);
  mapmech_xyconv_g520 : IND2D1BWP7T port map(A1 => lethaltile_y(3), B1 => lethaltile_y(0), ZN => mapmech_xyconv_n_3);
  mapmech_xyconv_g521 : INVD1BWP7T port map(I => lethaltile_x(1), ZN => mapmech_xyconv_n_2);
  mapmech_xyconv_g522 : INVD1BWP7T port map(I => lethaltile_y(1), ZN => mapmech_xyconv_n_1);
  mapmech_t38_g136 : BUFFD4BWP7T port map(I => mapmech_t38_state(1), Z => maptoVGA(166));
  mapmech_t38_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t38_n_7, A2 => mapmech_t38_n_8, Z => maptoVGA(167));
  mapmech_t38_g185 : NR2XD0BWP7T port map(A1 => mapmech_t38_n_4, A2 => n_0, ZN => mapmech_t38_n_6);
  mapmech_t38_g186 : AOI21D0BWP7T port map(A1 => mapmech_t38_n_2, A2 => mapmech_t38_n_3, B => n_0, ZN => mapmech_t38_n_5);
  mapmech_t38_g187 : AOI22D0BWP7T port map(A1 => mapmech_t38_state(1), A2 => mapmech_t38_n_3, B1 => mapmech_t38_state(0), B2 => mapmech_t38_n_1, ZN => mapmech_t38_n_4);
  mapmech_t38_g188 : ND3D0BWP7T port map(A1 => mapmech_yo3, A2 => mapmech_xo4, A3 => n_105, ZN => mapmech_t38_n_3);
  mapmech_t38_g189 : ND2D1BWP7T port map(A1 => mapmech_t38_state(0), A2 => n_105, ZN => mapmech_t38_n_2);
  mapmech_t38_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t38_n_1);
  mapmech_t38_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t38_n_5, Q => mapmech_t38_state(0), QN => mapmech_t38_n_8);
  mapmech_t38_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t38_n_6, Q => mapmech_t38_state(1), QN => mapmech_t38_n_7);
  mapmech_t39_g136 : BUFFD4BWP7T port map(I => mapmech_t39_state(1), Z => maptoVGA(164));
  mapmech_t39_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t39_n_7, A2 => mapmech_t39_n_9, Z => maptoVGA(165));
  mapmech_t39_g185 : NR2XD0BWP7T port map(A1 => mapmech_t39_n_4, A2 => n_0, ZN => mapmech_t39_n_6);
  mapmech_t39_g186 : AOI21D0BWP7T port map(A1 => mapmech_t39_n_2, A2 => mapmech_t39_n_3, B => n_0, ZN => mapmech_t39_n_5);
  mapmech_t39_g187 : AOI22D0BWP7T port map(A1 => mapmech_t39_state(1), A2 => mapmech_t39_n_3, B1 => mapmech_t39_state(0), B2 => mapmech_t39_n_1, ZN => mapmech_t39_n_4);
  mapmech_t39_g188 : ND3D0BWP7T port map(A1 => mapmech_xo5, A2 => mapmech_yo3, A3 => n_105, ZN => mapmech_t39_n_3);
  mapmech_t39_g189 : ND2D1BWP7T port map(A1 => mapmech_t39_state(0), A2 => n_105, ZN => mapmech_t39_n_2);
  mapmech_t39_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t39_n_1);
  mapmech_t39_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t39_n_5, Q => mapmech_t39_state(0), QN => mapmech_t39_n_9);
  mapmech_t39_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t39_n_6, Q => mapmech_t39_state(1), QN => mapmech_t39_n_7);
  mapmech_t40_g136 : BUFFD4BWP7T port map(I => mapmech_t40_state(1), Z => maptoVGA(162));
  mapmech_t40_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t40_n_7, A2 => mapmech_t40_n_8, Z => maptoVGA(163));
  mapmech_t40_g185 : NR2XD0BWP7T port map(A1 => mapmech_t40_n_4, A2 => n_0, ZN => mapmech_t40_n_6);
  mapmech_t40_g186 : AOI21D0BWP7T port map(A1 => mapmech_t40_n_2, A2 => mapmech_t40_n_3, B => n_0, ZN => mapmech_t40_n_5);
  mapmech_t40_g187 : AOI22D0BWP7T port map(A1 => mapmech_t40_state(1), A2 => mapmech_t40_n_3, B1 => mapmech_t40_state(0), B2 => mapmech_t40_n_1, ZN => mapmech_t40_n_4);
  mapmech_t40_g188 : ND3D0BWP7T port map(A1 => mapmech_yo3, A2 => mapmech_xo6, A3 => n_105, ZN => mapmech_t40_n_3);
  mapmech_t40_g189 : ND2D1BWP7T port map(A1 => mapmech_t40_state(0), A2 => n_105, ZN => mapmech_t40_n_2);
  mapmech_t40_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t40_n_1);
  mapmech_t40_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t40_n_5, Q => mapmech_t40_state(0), QN => mapmech_t40_n_8);
  mapmech_t40_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t40_n_6, Q => mapmech_t40_state(1), QN => mapmech_t40_n_7);
  mapmech_t41_g136 : BUFFD4BWP7T port map(I => mapmech_t41_state(1), Z => maptoVGA(160));
  mapmech_t41_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t41_n_7, A2 => mapmech_t41_n_8, Z => maptoVGA(161));
  mapmech_t41_g185 : NR2XD0BWP7T port map(A1 => mapmech_t41_n_4, A2 => n_0, ZN => mapmech_t41_n_6);
  mapmech_t41_g186 : AOI21D0BWP7T port map(A1 => mapmech_t41_n_2, A2 => mapmech_t41_n_3, B => n_0, ZN => mapmech_t41_n_5);
  mapmech_t41_g187 : AOI22D0BWP7T port map(A1 => mapmech_t41_state(1), A2 => mapmech_t41_n_3, B1 => mapmech_t41_state(0), B2 => mapmech_t41_n_1, ZN => mapmech_t41_n_4);
  mapmech_t41_g188 : ND3D0BWP7T port map(A1 => mapmech_xo7, A2 => mapmech_yo3, A3 => n_105, ZN => mapmech_t41_n_3);
  mapmech_t41_g189 : ND2D1BWP7T port map(A1 => mapmech_t41_state(0), A2 => n_105, ZN => mapmech_t41_n_2);
  mapmech_t41_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t41_n_1);
  mapmech_t41_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t41_n_5, Q => mapmech_t41_state(0), QN => mapmech_t41_n_8);
  mapmech_t41_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t41_n_6, Q => mapmech_t41_state(1), QN => mapmech_t41_n_7);
  mapmech_t42_g135 : BUFFD4BWP7T port map(I => mapmech_t42_state(1), Z => maptoVGA(158));
  mapmech_t42_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t42_n_7, A2 => mapmech_t42_n_8, Z => maptoVGA(159));
  mapmech_t42_g185 : NR2XD0BWP7T port map(A1 => mapmech_t42_n_4, A2 => n_0, ZN => mapmech_t42_n_6);
  mapmech_t42_g186 : AOI21D0BWP7T port map(A1 => mapmech_t42_n_2, A2 => mapmech_t42_n_3, B => n_0, ZN => mapmech_t42_n_5);
  mapmech_t42_g187 : AOI22D0BWP7T port map(A1 => mapmech_t42_state(1), A2 => mapmech_t42_n_3, B1 => mapmech_t42_state(0), B2 => mapmech_t42_n_1, ZN => mapmech_t42_n_4);
  mapmech_t42_g188 : ND3D0BWP7T port map(A1 => mapmech_yo3, A2 => mapmech_xo8, A3 => n_105, ZN => mapmech_t42_n_3);
  mapmech_t42_g189 : ND2D1BWP7T port map(A1 => mapmech_t42_state(0), A2 => n_105, ZN => mapmech_t42_n_2);
  mapmech_t42_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t42_n_1);
  mapmech_t42_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t42_n_5, Q => mapmech_t42_state(0), QN => mapmech_t42_n_8);
  mapmech_t42_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t42_n_6, Q => mapmech_t42_state(1), QN => mapmech_t42_n_7);
  mapmech_t43_g68 : INVD4BWP7T port map(I => mapmech_t43_state, ZN => maptoVGA(156));
  mapmech_t43_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t43_n_2, Q => mapmech_t43_state);
  mapmech_t43_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(156), A2 => mapmech_t43_n_1, B => n_0, C => mapmech_t43_n_0, ZN => mapmech_t43_n_2);
  mapmech_t43_g119 : ND2D0BWP7T port map(A1 => mapmech_yo3, A2 => mapmech_xo9, ZN => mapmech_t43_n_1);
  mapmech_t43_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t43_n_0);
  mapmech_t46_g135 : BUFFD4BWP7T port map(I => mapmech_t46_state(1), Z => maptoVGA(150));
  mapmech_t46_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t46_n_7, A2 => mapmech_t46_n_9, Z => maptoVGA(151));
  mapmech_t46_g185 : NR2XD0BWP7T port map(A1 => mapmech_t46_n_4, A2 => n_0, ZN => mapmech_t46_n_6);
  mapmech_t46_g186 : AOI21D0BWP7T port map(A1 => mapmech_t46_n_2, A2 => mapmech_t46_n_3, B => n_0, ZN => mapmech_t46_n_5);
  mapmech_t46_g187 : AOI22D0BWP7T port map(A1 => mapmech_t46_state(1), A2 => mapmech_t46_n_3, B1 => mapmech_t46_state(0), B2 => mapmech_t46_n_1, ZN => mapmech_t46_n_4);
  mapmech_t46_g188 : ND3D0BWP7T port map(A1 => mapmech_yo4, A2 => mapmech_xo1, A3 => n_105, ZN => mapmech_t46_n_3);
  mapmech_t46_g189 : ND2D1BWP7T port map(A1 => mapmech_t46_state(0), A2 => n_105, ZN => mapmech_t46_n_2);
  mapmech_t46_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t46_n_1);
  mapmech_t46_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t46_n_5, Q => mapmech_t46_state(0), QN => mapmech_t46_n_9);
  mapmech_t46_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t46_n_6, Q => mapmech_t46_state(1), QN => mapmech_t46_n_7);
  mapmech_t48_g136 : BUFFD4BWP7T port map(I => mapmech_t48_state(1), Z => maptoVGA(146));
  mapmech_t48_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t48_n_7, A2 => mapmech_t48_n_9, Z => maptoVGA(147));
  mapmech_t48_g185 : NR2XD0BWP7T port map(A1 => mapmech_t48_n_4, A2 => n_0, ZN => mapmech_t48_n_6);
  mapmech_t48_g186 : AOI21D0BWP7T port map(A1 => mapmech_t48_n_2, A2 => mapmech_t48_n_3, B => n_0, ZN => mapmech_t48_n_5);
  mapmech_t48_g187 : AOI22D0BWP7T port map(A1 => mapmech_t48_state(1), A2 => mapmech_t48_n_3, B1 => mapmech_t48_state(0), B2 => mapmech_t48_n_1, ZN => mapmech_t48_n_4);
  mapmech_t48_g188 : ND3D0BWP7T port map(A1 => mapmech_xo3, A2 => mapmech_yo4, A3 => n_105, ZN => mapmech_t48_n_3);
  mapmech_t48_g189 : ND2D1BWP7T port map(A1 => mapmech_t48_state(0), A2 => n_105, ZN => mapmech_t48_n_2);
  mapmech_t48_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t48_n_1);
  mapmech_t48_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t48_n_5, Q => mapmech_t48_state(0), QN => mapmech_t48_n_9);
  mapmech_t48_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t48_n_6, Q => mapmech_t48_state(1), QN => mapmech_t48_n_7);
  mapmech_t50_g68 : INVD4BWP7T port map(I => mapmech_t50_state, ZN => maptoVGA(142));
  mapmech_t50_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t50_n_2, Q => mapmech_t50_state);
  mapmech_t50_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(142), A2 => mapmech_t50_n_1, B => n_0, C => mapmech_t50_n_0, ZN => mapmech_t50_n_2);
  mapmech_t50_g119 : ND2D0BWP7T port map(A1 => mapmech_xo5, A2 => mapmech_yo4, ZN => mapmech_t50_n_1);
  mapmech_t50_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t50_n_0);
  mapmech_t52_g136 : BUFFD4BWP7T port map(I => mapmech_t52_state(1), Z => maptoVGA(138));
  mapmech_t52_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t52_n_7, A2 => mapmech_t52_n_9, Z => maptoVGA(139));
  mapmech_t52_g185 : NR2XD0BWP7T port map(A1 => mapmech_t52_n_4, A2 => n_0, ZN => mapmech_t52_n_6);
  mapmech_t52_g186 : AOI21D0BWP7T port map(A1 => mapmech_t52_n_2, A2 => mapmech_t52_n_3, B => n_0, ZN => mapmech_t52_n_5);
  mapmech_t52_g187 : AOI22D0BWP7T port map(A1 => mapmech_t52_state(1), A2 => mapmech_t52_n_3, B1 => mapmech_t52_state(0), B2 => mapmech_t52_n_1, ZN => mapmech_t52_n_4);
  mapmech_t52_g188 : ND3D0BWP7T port map(A1 => mapmech_xo7, A2 => mapmech_yo4, A3 => n_105, ZN => mapmech_t52_n_3);
  mapmech_t52_g189 : ND2D1BWP7T port map(A1 => mapmech_t52_state(0), A2 => n_105, ZN => mapmech_t52_n_2);
  mapmech_t52_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t52_n_1);
  mapmech_t52_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t52_n_5, Q => mapmech_t52_state(0), QN => mapmech_t52_n_9);
  mapmech_t52_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t52_n_6, Q => mapmech_t52_state(1), QN => mapmech_t52_n_7);
  mapmech_t54_g135 : BUFFD4BWP7T port map(I => mapmech_t54_state(1), Z => maptoVGA(134));
  mapmech_t54_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t54_n_7, A2 => mapmech_t54_n_8, Z => maptoVGA(135));
  mapmech_t54_g185 : NR2XD0BWP7T port map(A1 => mapmech_t54_n_4, A2 => n_0, ZN => mapmech_t54_n_6);
  mapmech_t54_g186 : AOI21D0BWP7T port map(A1 => mapmech_t54_n_2, A2 => mapmech_t54_n_3, B => n_0, ZN => mapmech_t54_n_5);
  mapmech_t54_g187 : AOI22D0BWP7T port map(A1 => mapmech_t54_state(1), A2 => mapmech_t54_n_3, B1 => mapmech_t54_state(0), B2 => mapmech_t54_n_1, ZN => mapmech_t54_n_4);
  mapmech_t54_g188 : ND3D0BWP7T port map(A1 => mapmech_yo4, A2 => mapmech_xo9, A3 => n_105, ZN => mapmech_t54_n_3);
  mapmech_t54_g189 : ND2D1BWP7T port map(A1 => mapmech_t54_state(0), A2 => n_105, ZN => mapmech_t54_n_2);
  mapmech_t54_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t54_n_1);
  mapmech_t54_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t54_n_5, Q => mapmech_t54_state(0), QN => mapmech_t54_n_8);
  mapmech_t54_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t54_n_6, Q => mapmech_t54_state(1), QN => mapmech_t54_n_7);
  mapmech_t57_g135 : BUFFD4BWP7T port map(I => mapmech_t57_state(1), Z => maptoVGA(128));
  mapmech_t57_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t57_n_7, A2 => mapmech_t57_n_9, Z => maptoVGA(129));
  mapmech_t57_g185 : NR2XD0BWP7T port map(A1 => mapmech_t57_n_4, A2 => n_0, ZN => mapmech_t57_n_6);
  mapmech_t57_g186 : AOI21D0BWP7T port map(A1 => mapmech_t57_n_2, A2 => mapmech_t57_n_3, B => n_0, ZN => mapmech_t57_n_5);
  mapmech_t57_g187 : AOI22D0BWP7T port map(A1 => mapmech_t57_state(1), A2 => mapmech_t57_n_3, B1 => mapmech_t57_state(0), B2 => mapmech_t57_n_1, ZN => mapmech_t57_n_4);
  mapmech_t57_g188 : ND3D0BWP7T port map(A1 => mapmech_yo5, A2 => mapmech_xo1, A3 => n_105, ZN => mapmech_t57_n_3);
  mapmech_t57_g189 : ND2D1BWP7T port map(A1 => mapmech_t57_state(0), A2 => n_105, ZN => mapmech_t57_n_2);
  mapmech_t57_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t57_n_1);
  mapmech_t57_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t57_n_5, Q => mapmech_t57_state(0), QN => mapmech_t57_n_9);
  mapmech_t57_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t57_n_6, Q => mapmech_t57_state(1), QN => mapmech_t57_n_7);
  mapmech_t58_g136 : BUFFD4BWP7T port map(I => mapmech_t58_state(1), Z => maptoVGA(126));
  mapmech_t58_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t58_n_7, A2 => mapmech_t58_n_8, Z => maptoVGA(127));
  mapmech_t58_g185 : NR2XD0BWP7T port map(A1 => mapmech_t58_n_4, A2 => n_0, ZN => mapmech_t58_n_6);
  mapmech_t58_g186 : AOI21D0BWP7T port map(A1 => mapmech_t58_n_2, A2 => mapmech_t58_n_3, B => n_0, ZN => mapmech_t58_n_5);
  mapmech_t58_g187 : AOI22D0BWP7T port map(A1 => mapmech_t58_state(1), A2 => mapmech_t58_n_3, B1 => mapmech_t58_state(0), B2 => mapmech_t58_n_1, ZN => mapmech_t58_n_4);
  mapmech_t58_g188 : ND3D0BWP7T port map(A1 => mapmech_yo5, A2 => mapmech_xo2, A3 => n_105, ZN => mapmech_t58_n_3);
  mapmech_t58_g189 : ND2D1BWP7T port map(A1 => mapmech_t58_state(0), A2 => n_105, ZN => mapmech_t58_n_2);
  mapmech_t58_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t58_n_1);
  mapmech_t58_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t58_n_5, Q => mapmech_t58_state(0), QN => mapmech_t58_n_8);
  mapmech_t58_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t58_n_6, Q => mapmech_t58_state(1), QN => mapmech_t58_n_7);
  mapmech_t59_g136 : BUFFD4BWP7T port map(I => mapmech_t59_state(1), Z => maptoVGA(124));
  mapmech_t59_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t59_n_7, A2 => mapmech_t59_n_8, Z => maptoVGA(125));
  mapmech_t59_g185 : NR2XD0BWP7T port map(A1 => mapmech_t59_n_4, A2 => n_0, ZN => mapmech_t59_n_6);
  mapmech_t59_g186 : AOI21D0BWP7T port map(A1 => mapmech_t59_n_2, A2 => mapmech_t59_n_3, B => n_0, ZN => mapmech_t59_n_5);
  mapmech_t59_g187 : AOI22D0BWP7T port map(A1 => mapmech_t59_state(1), A2 => mapmech_t59_n_3, B1 => mapmech_t59_state(0), B2 => mapmech_t59_n_1, ZN => mapmech_t59_n_4);
  mapmech_t59_g188 : ND3D0BWP7T port map(A1 => mapmech_yo5, A2 => mapmech_xo3, A3 => n_105, ZN => mapmech_t59_n_3);
  mapmech_t59_g189 : ND2D1BWP7T port map(A1 => mapmech_t59_state(0), A2 => n_105, ZN => mapmech_t59_n_2);
  mapmech_t59_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t59_n_1);
  mapmech_t59_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t59_n_5, Q => mapmech_t59_state(0), QN => mapmech_t59_n_8);
  mapmech_t59_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t59_n_6, Q => mapmech_t59_state(1), QN => mapmech_t59_n_7);
  mapmech_t60_g68 : INVD4BWP7T port map(I => mapmech_t60_state, ZN => maptoVGA(122));
  mapmech_t60_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t60_n_2, Q => mapmech_t60_state);
  mapmech_t60_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(122), A2 => mapmech_t60_n_1, B => n_0, C => mapmech_t60_n_0, ZN => mapmech_t60_n_2);
  mapmech_t60_g119 : ND2D0BWP7T port map(A1 => mapmech_yo5, A2 => mapmech_xo4, ZN => mapmech_t60_n_1);
  mapmech_t60_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t60_n_0);
  mapmech_t61_g68 : INVD4BWP7T port map(I => mapmech_t61_state, ZN => maptoVGA(120));
  mapmech_t61_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t61_n_2, Q => mapmech_t61_state);
  mapmech_t61_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(120), A2 => mapmech_t61_n_1, B => n_0, C => mapmech_t61_n_0, ZN => mapmech_t61_n_2);
  mapmech_t61_g119 : ND2D0BWP7T port map(A1 => mapmech_xo5, A2 => mapmech_yo5, ZN => mapmech_t61_n_1);
  mapmech_t61_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t61_n_0);
  mapmech_t62_g68 : INVD4BWP7T port map(I => mapmech_t62_state, ZN => maptoVGA(118));
  mapmech_t62_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t62_n_2, Q => mapmech_t62_state);
  mapmech_t62_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(118), A2 => mapmech_t62_n_1, B => n_0, C => mapmech_t62_n_0, ZN => mapmech_t62_n_2);
  mapmech_t62_g119 : ND2D0BWP7T port map(A1 => mapmech_yo5, A2 => mapmech_xo6, ZN => mapmech_t62_n_1);
  mapmech_t62_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t62_n_0);
  mapmech_t63_g136 : BUFFD4BWP7T port map(I => mapmech_t63_state(1), Z => maptoVGA(116));
  mapmech_t63_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t63_n_7, A2 => mapmech_t63_n_9, Z => maptoVGA(117));
  mapmech_t63_g185 : NR2XD0BWP7T port map(A1 => mapmech_t63_n_4, A2 => n_0, ZN => mapmech_t63_n_6);
  mapmech_t63_g186 : AOI21D0BWP7T port map(A1 => mapmech_t63_n_2, A2 => mapmech_t63_n_3, B => n_0, ZN => mapmech_t63_n_5);
  mapmech_t63_g187 : AOI22D0BWP7T port map(A1 => mapmech_t63_state(1), A2 => mapmech_t63_n_3, B1 => mapmech_t63_state(0), B2 => mapmech_t63_n_1, ZN => mapmech_t63_n_4);
  mapmech_t63_g188 : ND3D0BWP7T port map(A1 => mapmech_xo7, A2 => mapmech_yo5, A3 => n_105, ZN => mapmech_t63_n_3);
  mapmech_t63_g189 : ND2D1BWP7T port map(A1 => mapmech_t63_state(0), A2 => n_105, ZN => mapmech_t63_n_2);
  mapmech_t63_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t63_n_1);
  mapmech_t63_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t63_n_5, Q => mapmech_t63_state(0), QN => mapmech_t63_n_9);
  mapmech_t63_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t63_n_6, Q => mapmech_t63_state(1), QN => mapmech_t63_n_7);
  mapmech_t101_g68 : INVD4BWP7T port map(I => mapmech_t101_state, ZN => maptoVGA(40));
  mapmech_t101_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t101_n_2, Q => mapmech_t101_state);
  mapmech_t101_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(40), A2 => mapmech_t101_n_1, B => n_0, C => mapmech_t101_n_0, ZN => mapmech_t101_n_2);
  mapmech_t101_g119 : ND2D0BWP7T port map(A1 => mapmech_yo9, A2 => mapmech_xo1, ZN => mapmech_t101_n_1);
  mapmech_t101_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t101_n_0);
  mapmech_t64_g136 : BUFFD4BWP7T port map(I => mapmech_t64_state(1), Z => maptoVGA(114));
  mapmech_t64_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t64_n_7, A2 => mapmech_t64_n_9, Z => maptoVGA(115));
  mapmech_t64_g185 : NR2XD0BWP7T port map(A1 => mapmech_t64_n_4, A2 => n_0, ZN => mapmech_t64_n_6);
  mapmech_t64_g186 : AOI21D0BWP7T port map(A1 => mapmech_t64_n_2, A2 => mapmech_t64_n_3, B => n_0, ZN => mapmech_t64_n_5);
  mapmech_t64_g187 : AOI22D0BWP7T port map(A1 => mapmech_t64_state(1), A2 => mapmech_t64_n_3, B1 => mapmech_t64_state(0), B2 => mapmech_t64_n_1, ZN => mapmech_t64_n_4);
  mapmech_t64_g188 : ND3D0BWP7T port map(A1 => mapmech_yo5, A2 => mapmech_xo8, A3 => n_105, ZN => mapmech_t64_n_3);
  mapmech_t64_g189 : ND2D1BWP7T port map(A1 => mapmech_t64_state(0), A2 => n_105, ZN => mapmech_t64_n_2);
  mapmech_t64_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t64_n_1);
  mapmech_t64_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t64_n_5, Q => mapmech_t64_state(0), QN => mapmech_t64_n_9);
  mapmech_t64_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t64_n_6, Q => mapmech_t64_state(1), QN => mapmech_t64_n_7);
  mapmech_t102_g68 : INVD4BWP7T port map(I => mapmech_t102_state, ZN => maptoVGA(38));
  mapmech_t102_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t102_n_2, Q => mapmech_t102_state);
  mapmech_t102_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(38), A2 => mapmech_t102_n_1, B => n_0, C => mapmech_t102_n_0, ZN => mapmech_t102_n_2);
  mapmech_t102_g119 : ND2D0BWP7T port map(A1 => mapmech_yo9, A2 => mapmech_xo2, ZN => mapmech_t102_n_1);
  mapmech_t102_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t102_n_0);
  mapmech_t65_g136 : BUFFD4BWP7T port map(I => mapmech_t65_state(1), Z => maptoVGA(112));
  mapmech_t65_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t65_n_7, A2 => mapmech_t65_n_9, Z => maptoVGA(113));
  mapmech_t65_g185 : NR2XD0BWP7T port map(A1 => mapmech_t65_n_4, A2 => n_0, ZN => mapmech_t65_n_6);
  mapmech_t65_g186 : AOI21D0BWP7T port map(A1 => mapmech_t65_n_2, A2 => mapmech_t65_n_3, B => n_0, ZN => mapmech_t65_n_5);
  mapmech_t65_g187 : AOI22D0BWP7T port map(A1 => mapmech_t65_state(1), A2 => mapmech_t65_n_3, B1 => mapmech_t65_state(0), B2 => mapmech_t65_n_1, ZN => mapmech_t65_n_4);
  mapmech_t65_g188 : ND3D0BWP7T port map(A1 => mapmech_yo5, A2 => mapmech_xo9, A3 => n_105, ZN => mapmech_t65_n_3);
  mapmech_t65_g189 : ND2D1BWP7T port map(A1 => mapmech_t65_state(0), A2 => n_105, ZN => mapmech_t65_n_2);
  mapmech_t65_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t65_n_1);
  mapmech_t65_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t65_n_5, Q => mapmech_t65_state(0), QN => mapmech_t65_n_9);
  mapmech_t65_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t65_n_6, Q => mapmech_t65_state(1), QN => mapmech_t65_n_7);
  mapmech_t103_g68 : INVD4BWP7T port map(I => mapmech_t103_state, ZN => maptoVGA(36));
  mapmech_t103_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t103_n_2, Q => mapmech_t103_state);
  mapmech_t103_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(36), A2 => mapmech_t103_n_1, B => n_0, C => mapmech_t103_n_0, ZN => mapmech_t103_n_2);
  mapmech_t103_g119 : ND2D0BWP7T port map(A1 => mapmech_xo3, A2 => mapmech_yo9, ZN => mapmech_t103_n_1);
  mapmech_t103_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t103_n_0);
  mapmech_t104_g136 : BUFFD4BWP7T port map(I => mapmech_t104_state(1), Z => maptoVGA(34));
  mapmech_t104_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t104_n_7, A2 => mapmech_t104_n_9, Z => maptoVGA(35));
  mapmech_t104_g185 : NR2XD0BWP7T port map(A1 => mapmech_t104_n_4, A2 => n_0, ZN => mapmech_t104_n_6);
  mapmech_t104_g186 : AOI21D0BWP7T port map(A1 => mapmech_t104_n_2, A2 => mapmech_t104_n_3, B => n_0, ZN => mapmech_t104_n_5);
  mapmech_t104_g187 : AOI22D0BWP7T port map(A1 => mapmech_t104_state(1), A2 => mapmech_t104_n_3, B1 => mapmech_t104_state(0), B2 => mapmech_t104_n_1, ZN => mapmech_t104_n_4);
  mapmech_t104_g188 : ND3D0BWP7T port map(A1 => mapmech_xo4, A2 => mapmech_yo9, A3 => n_105, ZN => mapmech_t104_n_3);
  mapmech_t104_g189 : ND2D1BWP7T port map(A1 => mapmech_t104_state(0), A2 => n_105, ZN => mapmech_t104_n_2);
  mapmech_t104_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t104_n_1);
  mapmech_t104_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t104_n_5, Q => mapmech_t104_state(0), QN => mapmech_t104_n_9);
  mapmech_t104_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t104_n_6, Q => mapmech_t104_state(1), QN => mapmech_t104_n_7);
  mapmech_t105_g136 : BUFFD4BWP7T port map(I => mapmech_t105_state(1), Z => maptoVGA(32));
  mapmech_t105_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t105_n_7, A2 => mapmech_t105_n_9, Z => maptoVGA(33));
  mapmech_t105_g185 : NR2XD0BWP7T port map(A1 => mapmech_t105_n_4, A2 => n_0, ZN => mapmech_t105_n_6);
  mapmech_t105_g186 : AOI21D0BWP7T port map(A1 => mapmech_t105_n_2, A2 => mapmech_t105_n_3, B => n_0, ZN => mapmech_t105_n_5);
  mapmech_t105_g187 : AOI22D0BWP7T port map(A1 => mapmech_t105_state(1), A2 => mapmech_t105_n_3, B1 => mapmech_t105_state(0), B2 => mapmech_t105_n_1, ZN => mapmech_t105_n_4);
  mapmech_t105_g188 : ND3D0BWP7T port map(A1 => mapmech_xo5, A2 => mapmech_yo9, A3 => n_105, ZN => mapmech_t105_n_3);
  mapmech_t105_g189 : ND2D1BWP7T port map(A1 => mapmech_t105_state(0), A2 => n_105, ZN => mapmech_t105_n_2);
  mapmech_t105_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t105_n_1);
  mapmech_t105_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t105_n_5, Q => mapmech_t105_state(0), QN => mapmech_t105_n_9);
  mapmech_t105_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t105_n_6, Q => mapmech_t105_state(1), QN => mapmech_t105_n_7);
  mapmech_t68_g136 : BUFFD4BWP7T port map(I => mapmech_t68_state(1), Z => maptoVGA(106));
  mapmech_t68_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t68_n_7, A2 => mapmech_t68_n_8, Z => maptoVGA(107));
  mapmech_t68_g185 : NR2XD0BWP7T port map(A1 => mapmech_t68_n_4, A2 => n_0, ZN => mapmech_t68_n_6);
  mapmech_t68_g186 : AOI21D0BWP7T port map(A1 => mapmech_t68_n_2, A2 => mapmech_t68_n_3, B => n_0, ZN => mapmech_t68_n_5);
  mapmech_t68_g187 : AOI22D0BWP7T port map(A1 => mapmech_t68_state(1), A2 => mapmech_t68_n_3, B1 => mapmech_t68_state(0), B2 => mapmech_t68_n_1, ZN => mapmech_t68_n_4);
  mapmech_t68_g188 : ND3D0BWP7T port map(A1 => mapmech_yo6, A2 => mapmech_xo1, A3 => n_105, ZN => mapmech_t68_n_3);
  mapmech_t68_g189 : ND2D1BWP7T port map(A1 => mapmech_t68_state(0), A2 => n_105, ZN => mapmech_t68_n_2);
  mapmech_t68_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t68_n_1);
  mapmech_t68_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t68_n_5, Q => mapmech_t68_state(0), QN => mapmech_t68_n_8);
  mapmech_t68_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t68_n_6, Q => mapmech_t68_state(1), QN => mapmech_t68_n_7);
  mapmech_t106_g136 : BUFFD4BWP7T port map(I => mapmech_t106_state(1), Z => maptoVGA(30));
  mapmech_t106_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t106_n_7, A2 => mapmech_t106_n_8, Z => maptoVGA(31));
  mapmech_t106_g185 : NR2XD0BWP7T port map(A1 => mapmech_t106_n_4, A2 => n_0, ZN => mapmech_t106_n_6);
  mapmech_t106_g186 : AOI21D0BWP7T port map(A1 => mapmech_t106_n_2, A2 => mapmech_t106_n_3, B => n_0, ZN => mapmech_t106_n_5);
  mapmech_t106_g187 : AOI22D0BWP7T port map(A1 => mapmech_t106_state(1), A2 => mapmech_t106_n_3, B1 => mapmech_t106_state(0), B2 => mapmech_t106_n_1, ZN => mapmech_t106_n_4);
  mapmech_t106_g188 : ND3D0BWP7T port map(A1 => mapmech_xo6, A2 => mapmech_yo9, A3 => n_105, ZN => mapmech_t106_n_3);
  mapmech_t106_g189 : ND2D1BWP7T port map(A1 => mapmech_t106_state(0), A2 => n_105, ZN => mapmech_t106_n_2);
  mapmech_t106_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t106_n_1);
  mapmech_t106_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t106_n_5, Q => mapmech_t106_state(0), QN => mapmech_t106_n_8);
  mapmech_t106_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t106_n_6, Q => mapmech_t106_state(1), QN => mapmech_t106_n_7);
  mapmech_t70_g136 : BUFFD4BWP7T port map(I => mapmech_t70_state(1), Z => maptoVGA(102));
  mapmech_t70_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t70_n_7, A2 => mapmech_t70_n_9, Z => maptoVGA(103));
  mapmech_t70_g185 : NR2XD0BWP7T port map(A1 => mapmech_t70_n_4, A2 => n_0, ZN => mapmech_t70_n_6);
  mapmech_t70_g186 : AOI21D0BWP7T port map(A1 => mapmech_t70_n_2, A2 => mapmech_t70_n_3, B => n_0, ZN => mapmech_t70_n_5);
  mapmech_t70_g187 : AOI22D0BWP7T port map(A1 => mapmech_t70_state(1), A2 => mapmech_t70_n_3, B1 => mapmech_t70_state(0), B2 => mapmech_t70_n_1, ZN => mapmech_t70_n_4);
  mapmech_t70_g188 : ND3D0BWP7T port map(A1 => mapmech_xo3, A2 => mapmech_yo6, A3 => n_105, ZN => mapmech_t70_n_3);
  mapmech_t70_g189 : ND2D1BWP7T port map(A1 => mapmech_t70_state(0), A2 => n_105, ZN => mapmech_t70_n_2);
  mapmech_t70_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t70_n_1);
  mapmech_t70_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t70_n_5, Q => mapmech_t70_state(0), QN => mapmech_t70_n_9);
  mapmech_t70_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t70_n_6, Q => mapmech_t70_state(1), QN => mapmech_t70_n_7);
  mapmech_t107_g68 : INVD4BWP7T port map(I => mapmech_t107_state, ZN => maptoVGA(28));
  mapmech_t107_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t107_n_2, Q => mapmech_t107_state);
  mapmech_t107_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(28), A2 => mapmech_t107_n_1, B => n_0, C => mapmech_t107_n_0, ZN => mapmech_t107_n_2);
  mapmech_t107_g119 : ND2D0BWP7T port map(A1 => mapmech_xo7, A2 => mapmech_yo9, ZN => mapmech_t107_n_1);
  mapmech_t107_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t107_n_0);
  mapmech_t108_g68 : INVD4BWP7T port map(I => mapmech_t108_state, ZN => maptoVGA(26));
  mapmech_t108_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t108_n_2, Q => mapmech_t108_state);
  mapmech_t108_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(26), A2 => mapmech_t108_n_1, B => n_0, C => mapmech_t108_n_0, ZN => mapmech_t108_n_2);
  mapmech_t108_g119 : ND2D0BWP7T port map(A1 => mapmech_yo9, A2 => mapmech_xo8, ZN => mapmech_t108_n_1);
  mapmech_t108_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t108_n_0);
  mapmech_t72_g68 : INVD4BWP7T port map(I => mapmech_t72_state, ZN => maptoVGA(98));
  mapmech_t72_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t72_n_2, Q => mapmech_t72_state);
  mapmech_t72_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(98), A2 => mapmech_t72_n_1, B => n_0, C => mapmech_t72_n_0, ZN => mapmech_t72_n_2);
  mapmech_t72_g119 : ND2D0BWP7T port map(A1 => mapmech_xo5, A2 => mapmech_yo6, ZN => mapmech_t72_n_1);
  mapmech_t72_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t72_n_0);
  mapmech_t109_g68 : INVD4BWP7T port map(I => mapmech_t109_state, ZN => maptoVGA(24));
  mapmech_t109_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t109_n_2, Q => mapmech_t109_state);
  mapmech_t109_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(24), A2 => mapmech_t109_n_1, B => n_0, C => mapmech_t109_n_0, ZN => mapmech_t109_n_2);
  mapmech_t109_g119 : ND2D0BWP7T port map(A1 => mapmech_yo9, A2 => mapmech_xo9, ZN => mapmech_t109_n_1);
  mapmech_t109_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t109_n_0);
  mapmech_t74_g136 : BUFFD4BWP7T port map(I => mapmech_t74_state(1), Z => maptoVGA(94));
  mapmech_t74_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t74_n_7, A2 => mapmech_t74_n_9, Z => maptoVGA(95));
  mapmech_t74_g185 : NR2XD0BWP7T port map(A1 => mapmech_t74_n_4, A2 => n_0, ZN => mapmech_t74_n_6);
  mapmech_t74_g186 : AOI21D0BWP7T port map(A1 => mapmech_t74_n_2, A2 => mapmech_t74_n_3, B => n_0, ZN => mapmech_t74_n_5);
  mapmech_t74_g187 : AOI22D0BWP7T port map(A1 => mapmech_t74_state(1), A2 => mapmech_t74_n_3, B1 => mapmech_t74_state(0), B2 => mapmech_t74_n_1, ZN => mapmech_t74_n_4);
  mapmech_t74_g188 : ND3D0BWP7T port map(A1 => mapmech_xo7, A2 => mapmech_yo6, A3 => n_105, ZN => mapmech_t74_n_3);
  mapmech_t74_g189 : ND2D1BWP7T port map(A1 => mapmech_t74_state(0), A2 => n_105, ZN => mapmech_t74_n_2);
  mapmech_t74_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t74_n_1);
  mapmech_t74_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t74_n_5, Q => mapmech_t74_state(0), QN => mapmech_t74_n_9);
  mapmech_t74_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t74_n_6, Q => mapmech_t74_state(1), QN => mapmech_t74_n_7);
  mapmech_t76_g135 : BUFFD4BWP7T port map(I => mapmech_t76_state(1), Z => maptoVGA(90));
  mapmech_t76_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t76_n_7, A2 => mapmech_t76_n_9, Z => maptoVGA(91));
  mapmech_t76_g185 : NR2XD0BWP7T port map(A1 => mapmech_t76_n_4, A2 => n_0, ZN => mapmech_t76_n_6);
  mapmech_t76_g186 : AOI21D0BWP7T port map(A1 => mapmech_t76_n_2, A2 => mapmech_t76_n_3, B => n_0, ZN => mapmech_t76_n_5);
  mapmech_t76_g187 : AOI22D0BWP7T port map(A1 => mapmech_t76_state(1), A2 => mapmech_t76_n_3, B1 => mapmech_t76_state(0), B2 => mapmech_t76_n_1, ZN => mapmech_t76_n_4);
  mapmech_t76_g188 : ND3D0BWP7T port map(A1 => mapmech_yo6, A2 => mapmech_xo9, A3 => n_105, ZN => mapmech_t76_n_3);
  mapmech_t76_g189 : ND2D1BWP7T port map(A1 => mapmech_t76_state(0), A2 => n_105, ZN => mapmech_t76_n_2);
  mapmech_t76_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t76_n_1);
  mapmech_t76_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t76_n_5, Q => mapmech_t76_state(0), QN => mapmech_t76_n_9);
  mapmech_t76_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t76_n_6, Q => mapmech_t76_state(1), QN => mapmech_t76_n_7);
  mapmech_t80_g135 : BUFFD4BWP7T port map(I => mapmech_t80_state(1), Z => maptoVGA(82));
  mapmech_t80_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t80_n_7, A2 => mapmech_t80_n_9, Z => maptoVGA(83));
  mapmech_t80_g185 : NR2XD0BWP7T port map(A1 => mapmech_t80_n_4, A2 => n_0, ZN => mapmech_t80_n_6);
  mapmech_t80_g186 : AOI21D0BWP7T port map(A1 => mapmech_t80_n_2, A2 => mapmech_t80_n_3, B => n_0, ZN => mapmech_t80_n_5);
  mapmech_t80_g187 : AOI22D0BWP7T port map(A1 => mapmech_t80_state(1), A2 => mapmech_t80_n_3, B1 => mapmech_t80_state(0), B2 => mapmech_t80_n_1, ZN => mapmech_t80_n_4);
  mapmech_t80_g188 : ND3D0BWP7T port map(A1 => mapmech_yo7, A2 => mapmech_xo2, A3 => n_105, ZN => mapmech_t80_n_3);
  mapmech_t80_g189 : ND2D1BWP7T port map(A1 => mapmech_t80_state(0), A2 => n_105, ZN => mapmech_t80_n_2);
  mapmech_t80_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t80_n_1);
  mapmech_t80_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t80_n_5, Q => mapmech_t80_state(0), QN => mapmech_t80_n_9);
  mapmech_t80_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t80_n_6, Q => mapmech_t80_state(1), QN => mapmech_t80_n_7);
  mapmech_t79_g68 : INVD4BWP7T port map(I => mapmech_t79_state, ZN => maptoVGA(84));
  mapmech_t79_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t79_n_2, Q => mapmech_t79_state);
  mapmech_t79_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(84), A2 => mapmech_t79_n_1, B => n_0, C => mapmech_t79_n_0, ZN => mapmech_t79_n_2);
  mapmech_t79_g119 : ND2D0BWP7T port map(A1 => mapmech_yo7, A2 => mapmech_xo1, ZN => mapmech_t79_n_1);
  mapmech_t79_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t79_n_0);
  mapmech_t81_g135 : BUFFD4BWP7T port map(I => mapmech_t81_state(1), Z => maptoVGA(80));
  mapmech_t81_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t81_n_7, A2 => mapmech_t81_n_8, Z => maptoVGA(81));
  mapmech_t81_g185 : NR2XD0BWP7T port map(A1 => mapmech_t81_n_4, A2 => n_0, ZN => mapmech_t81_n_6);
  mapmech_t81_g186 : AOI21D0BWP7T port map(A1 => mapmech_t81_n_2, A2 => mapmech_t81_n_3, B => n_0, ZN => mapmech_t81_n_5);
  mapmech_t81_g187 : AOI22D0BWP7T port map(A1 => mapmech_t81_state(1), A2 => mapmech_t81_n_3, B1 => mapmech_t81_state(0), B2 => mapmech_t81_n_1, ZN => mapmech_t81_n_4);
  mapmech_t81_g188 : ND3D0BWP7T port map(A1 => mapmech_yo7, A2 => mapmech_xo3, A3 => n_105, ZN => mapmech_t81_n_3);
  mapmech_t81_g189 : ND2D1BWP7T port map(A1 => mapmech_t81_state(0), A2 => n_105, ZN => mapmech_t81_n_2);
  mapmech_t81_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t81_n_1);
  mapmech_t81_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t81_n_5, Q => mapmech_t81_state(0), QN => mapmech_t81_n_8);
  mapmech_t81_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t81_n_6, Q => mapmech_t81_state(1), QN => mapmech_t81_n_7);
  mapmech_t82_g136 : BUFFD4BWP7T port map(I => mapmech_t82_state(1), Z => maptoVGA(78));
  mapmech_t82_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t82_n_7, A2 => mapmech_t82_n_8, Z => maptoVGA(79));
  mapmech_t82_g185 : NR2XD0BWP7T port map(A1 => mapmech_t82_n_4, A2 => n_0, ZN => mapmech_t82_n_6);
  mapmech_t82_g186 : AOI21D0BWP7T port map(A1 => mapmech_t82_n_2, A2 => mapmech_t82_n_3, B => n_0, ZN => mapmech_t82_n_5);
  mapmech_t82_g187 : AOI22D0BWP7T port map(A1 => mapmech_t82_state(1), A2 => mapmech_t82_n_3, B1 => mapmech_t82_state(0), B2 => mapmech_t82_n_1, ZN => mapmech_t82_n_4);
  mapmech_t82_g188 : ND3D0BWP7T port map(A1 => mapmech_yo7, A2 => mapmech_xo4, A3 => n_105, ZN => mapmech_t82_n_3);
  mapmech_t82_g189 : ND2D1BWP7T port map(A1 => mapmech_t82_state(0), A2 => n_105, ZN => mapmech_t82_n_2);
  mapmech_t82_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t82_n_1);
  mapmech_t82_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t82_n_5, Q => mapmech_t82_state(0), QN => mapmech_t82_n_8);
  mapmech_t82_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t82_n_6, Q => mapmech_t82_state(1), QN => mapmech_t82_n_7);
  mapmech_t83_g136 : BUFFD4BWP7T port map(I => mapmech_t83_state(1), Z => maptoVGA(76));
  mapmech_t83_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t83_n_7, A2 => mapmech_t83_n_8, Z => maptoVGA(77));
  mapmech_t83_g185 : NR2XD0BWP7T port map(A1 => mapmech_t83_n_4, A2 => n_0, ZN => mapmech_t83_n_6);
  mapmech_t83_g186 : AOI21D0BWP7T port map(A1 => mapmech_t83_n_2, A2 => mapmech_t83_n_3, B => n_0, ZN => mapmech_t83_n_5);
  mapmech_t83_g187 : AOI22D0BWP7T port map(A1 => mapmech_t83_state(1), A2 => mapmech_t83_n_3, B1 => mapmech_t83_state(0), B2 => mapmech_t83_n_1, ZN => mapmech_t83_n_4);
  mapmech_t83_g188 : ND3D0BWP7T port map(A1 => mapmech_xo5, A2 => mapmech_yo7, A3 => n_105, ZN => mapmech_t83_n_3);
  mapmech_t83_g189 : ND2D1BWP7T port map(A1 => mapmech_t83_state(0), A2 => n_105, ZN => mapmech_t83_n_2);
  mapmech_t83_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t83_n_1);
  mapmech_t83_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t83_n_5, Q => mapmech_t83_state(0), QN => mapmech_t83_n_8);
  mapmech_t83_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t83_n_6, Q => mapmech_t83_state(1), QN => mapmech_t83_n_7);
  mapmech_t84_g136 : BUFFD4BWP7T port map(I => mapmech_t84_state(1), Z => maptoVGA(74));
  mapmech_t84_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t84_n_7, A2 => mapmech_t84_n_9, Z => maptoVGA(75));
  mapmech_t84_g185 : NR2XD0BWP7T port map(A1 => mapmech_t84_n_4, A2 => n_0, ZN => mapmech_t84_n_6);
  mapmech_t84_g186 : AOI21D0BWP7T port map(A1 => mapmech_t84_n_2, A2 => mapmech_t84_n_3, B => n_0, ZN => mapmech_t84_n_5);
  mapmech_t84_g187 : AOI22D0BWP7T port map(A1 => mapmech_t84_state(1), A2 => mapmech_t84_n_3, B1 => mapmech_t84_state(0), B2 => mapmech_t84_n_1, ZN => mapmech_t84_n_4);
  mapmech_t84_g188 : ND3D0BWP7T port map(A1 => mapmech_yo7, A2 => mapmech_xo6, A3 => n_105, ZN => mapmech_t84_n_3);
  mapmech_t84_g189 : ND2D1BWP7T port map(A1 => mapmech_t84_state(0), A2 => n_105, ZN => mapmech_t84_n_2);
  mapmech_t84_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t84_n_1);
  mapmech_t84_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t84_n_5, Q => mapmech_t84_state(0), QN => mapmech_t84_n_9);
  mapmech_t84_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t84_n_6, Q => mapmech_t84_state(1), QN => mapmech_t84_n_7);
  mapmech_t13_g68 : INVD4BWP7T port map(I => mapmech_t13_state, ZN => maptoVGA(216));
  mapmech_t13_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t13_n_2, Q => mapmech_t13_state);
  mapmech_t13_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(216), A2 => mapmech_t13_n_1, B => n_0, C => mapmech_t13_n_0, ZN => mapmech_t13_n_2);
  mapmech_t13_g119 : ND2D0BWP7T port map(A1 => mapmech_xo1, A2 => mapmech_yo1, ZN => mapmech_t13_n_1);
  mapmech_t13_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t13_n_0);
  mapmech_t85_g136 : BUFFD4BWP7T port map(I => mapmech_t85_state(1), Z => maptoVGA(72));
  mapmech_t85_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t85_n_7, A2 => mapmech_t85_n_9, Z => maptoVGA(73));
  mapmech_t85_g185 : NR2XD0BWP7T port map(A1 => mapmech_t85_n_4, A2 => n_0, ZN => mapmech_t85_n_6);
  mapmech_t85_g186 : AOI21D0BWP7T port map(A1 => mapmech_t85_n_2, A2 => mapmech_t85_n_3, B => n_0, ZN => mapmech_t85_n_5);
  mapmech_t85_g187 : AOI22D0BWP7T port map(A1 => mapmech_t85_state(1), A2 => mapmech_t85_n_3, B1 => mapmech_t85_state(0), B2 => mapmech_t85_n_1, ZN => mapmech_t85_n_4);
  mapmech_t85_g188 : ND3D0BWP7T port map(A1 => mapmech_xo7, A2 => mapmech_yo7, A3 => n_105, ZN => mapmech_t85_n_3);
  mapmech_t85_g189 : ND2D1BWP7T port map(A1 => mapmech_t85_state(0), A2 => n_105, ZN => mapmech_t85_n_2);
  mapmech_t85_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t85_n_1);
  mapmech_t85_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t85_n_5, Q => mapmech_t85_state(0), QN => mapmech_t85_n_9);
  mapmech_t85_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t85_n_6, Q => mapmech_t85_state(1), QN => mapmech_t85_n_7);
  mapmech_t14_g68 : INVD4BWP7T port map(I => mapmech_t14_state, ZN => maptoVGA(214));
  mapmech_t14_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t14_n_2, Q => mapmech_t14_state);
  mapmech_t14_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(214), A2 => mapmech_t14_n_1, B => n_0, C => mapmech_t14_n_0, ZN => mapmech_t14_n_2);
  mapmech_t14_g119 : ND2D0BWP7T port map(A1 => mapmech_yo1, A2 => mapmech_xo2, ZN => mapmech_t14_n_1);
  mapmech_t14_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t14_n_0);
  mapmech_t86_g136 : BUFFD4BWP7T port map(I => mapmech_t86_state(1), Z => maptoVGA(70));
  mapmech_t86_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t86_n_7, A2 => mapmech_t86_n_8, Z => maptoVGA(71));
  mapmech_t86_g185 : NR2XD0BWP7T port map(A1 => mapmech_t86_n_4, A2 => n_0, ZN => mapmech_t86_n_6);
  mapmech_t86_g186 : AOI21D0BWP7T port map(A1 => mapmech_t86_n_2, A2 => mapmech_t86_n_3, B => n_0, ZN => mapmech_t86_n_5);
  mapmech_t86_g187 : AOI22D0BWP7T port map(A1 => mapmech_t86_state(1), A2 => mapmech_t86_n_3, B1 => mapmech_t86_state(0), B2 => mapmech_t86_n_1, ZN => mapmech_t86_n_4);
  mapmech_t86_g188 : ND3D0BWP7T port map(A1 => mapmech_yo7, A2 => mapmech_xo8, A3 => n_105, ZN => mapmech_t86_n_3);
  mapmech_t86_g189 : ND2D1BWP7T port map(A1 => mapmech_t86_state(0), A2 => n_105, ZN => mapmech_t86_n_2);
  mapmech_t86_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t86_n_1);
  mapmech_t86_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t86_n_5, Q => mapmech_t86_state(0), QN => mapmech_t86_n_8);
  mapmech_t86_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t86_n_6, Q => mapmech_t86_state(1), QN => mapmech_t86_n_7);
  mapmech_t15_g68 : INVD4BWP7T port map(I => mapmech_t15_state, ZN => maptoVGA(212));
  mapmech_t15_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t15_n_2, Q => mapmech_t15_state);
  mapmech_t15_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(212), A2 => mapmech_t15_n_1, B => n_0, C => mapmech_t15_n_0, ZN => mapmech_t15_n_2);
  mapmech_t15_g119 : ND2D0BWP7T port map(A1 => mapmech_xo3, A2 => mapmech_yo1, ZN => mapmech_t15_n_1);
  mapmech_t15_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t15_n_0);
  mapmech_t87_g68 : INVD4BWP7T port map(I => mapmech_t87_state, ZN => maptoVGA(68));
  mapmech_t87_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t87_n_2, Q => mapmech_t87_state);
  mapmech_t87_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(68), A2 => mapmech_t87_n_1, B => n_0, C => mapmech_t87_n_0, ZN => mapmech_t87_n_2);
  mapmech_t87_g119 : ND2D0BWP7T port map(A1 => mapmech_yo7, A2 => mapmech_xo9, ZN => mapmech_t87_n_1);
  mapmech_t87_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t87_n_0);
  mapmech_t16_g136 : BUFFD4BWP7T port map(I => mapmech_t16_state(1), Z => maptoVGA(210));
  mapmech_t16_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t16_n_7, A2 => mapmech_t16_n_8, Z => maptoVGA(211));
  mapmech_t16_g185 : NR2XD0BWP7T port map(A1 => mapmech_t16_n_4, A2 => n_0, ZN => mapmech_t16_n_6);
  mapmech_t16_g186 : AOI21D0BWP7T port map(A1 => mapmech_t16_n_2, A2 => mapmech_t16_n_3, B => n_0, ZN => mapmech_t16_n_5);
  mapmech_t16_g187 : AOI22D0BWP7T port map(A1 => mapmech_t16_state(1), A2 => mapmech_t16_n_3, B1 => mapmech_t16_state(0), B2 => mapmech_t16_n_1, ZN => mapmech_t16_n_4);
  mapmech_t16_g188 : ND3D0BWP7T port map(A1 => mapmech_xo4, A2 => mapmech_yo1, A3 => n_105, ZN => mapmech_t16_n_3);
  mapmech_t16_g189 : ND2D1BWP7T port map(A1 => mapmech_t16_state(0), A2 => n_105, ZN => mapmech_t16_n_2);
  mapmech_t16_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t16_n_1);
  mapmech_t16_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t16_n_5, Q => mapmech_t16_state(0), QN => mapmech_t16_n_8);
  mapmech_t16_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t16_n_6, Q => mapmech_t16_state(1), QN => mapmech_t16_n_7);
  mapmech_t17_g135 : BUFFD4BWP7T port map(I => mapmech_t17_state(1), Z => maptoVGA(208));
  mapmech_t17_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t17_n_7, A2 => mapmech_t17_n_9, Z => maptoVGA(209));
  mapmech_t17_g185 : NR2XD0BWP7T port map(A1 => mapmech_t17_n_4, A2 => n_0, ZN => mapmech_t17_n_6);
  mapmech_t17_g186 : AOI21D0BWP7T port map(A1 => mapmech_t17_n_2, A2 => mapmech_t17_n_3, B => n_0, ZN => mapmech_t17_n_5);
  mapmech_t17_g187 : AOI22D0BWP7T port map(A1 => mapmech_t17_state(1), A2 => mapmech_t17_n_3, B1 => mapmech_t17_state(0), B2 => mapmech_t17_n_1, ZN => mapmech_t17_n_4);
  mapmech_t17_g188 : ND3D0BWP7T port map(A1 => mapmech_xo5, A2 => mapmech_yo1, A3 => n_105, ZN => mapmech_t17_n_3);
  mapmech_t17_g189 : ND2D1BWP7T port map(A1 => mapmech_t17_state(0), A2 => n_105, ZN => mapmech_t17_n_2);
  mapmech_t17_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t17_n_1);
  mapmech_t17_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t17_n_5, Q => mapmech_t17_state(0), QN => mapmech_t17_n_9);
  mapmech_t17_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t17_n_6, Q => mapmech_t17_state(1), QN => mapmech_t17_n_7);
  mapmech_t90_g68 : INVD4BWP7T port map(I => mapmech_t90_state, ZN => maptoVGA(62));
  mapmech_t90_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t90_n_2, Q => mapmech_t90_state);
  mapmech_t90_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(62), A2 => mapmech_t90_n_1, B => n_0, C => mapmech_t90_n_0, ZN => mapmech_t90_n_2);
  mapmech_t90_g119 : ND2D0BWP7T port map(A1 => mapmech_yo8, A2 => mapmech_xo1, ZN => mapmech_t90_n_1);
  mapmech_t90_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t90_n_0);
  mapmech_t18_g136 : BUFFD4BWP7T port map(I => mapmech_t18_state(1), Z => maptoVGA(206));
  mapmech_t18_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t18_n_7, A2 => mapmech_t18_n_8, Z => maptoVGA(207));
  mapmech_t18_g185 : NR2XD0BWP7T port map(A1 => mapmech_t18_n_4, A2 => n_0, ZN => mapmech_t18_n_6);
  mapmech_t18_g186 : AOI21D0BWP7T port map(A1 => mapmech_t18_n_2, A2 => mapmech_t18_n_3, B => n_0, ZN => mapmech_t18_n_5);
  mapmech_t18_g187 : AOI22D0BWP7T port map(A1 => mapmech_t18_state(1), A2 => mapmech_t18_n_3, B1 => mapmech_t18_state(0), B2 => mapmech_t18_n_1, ZN => mapmech_t18_n_4);
  mapmech_t18_g188 : ND3D0BWP7T port map(A1 => mapmech_xo6, A2 => mapmech_yo1, A3 => n_105, ZN => mapmech_t18_n_3);
  mapmech_t18_g189 : ND2D1BWP7T port map(A1 => mapmech_t18_state(0), A2 => n_105, ZN => mapmech_t18_n_2);
  mapmech_t18_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t18_n_1);
  mapmech_t18_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t18_n_5, Q => mapmech_t18_state(0), QN => mapmech_t18_n_8);
  mapmech_t18_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t18_n_6, Q => mapmech_t18_state(1), QN => mapmech_t18_n_7);
  mapmech_t19_g68 : INVD4BWP7T port map(I => mapmech_t19_state, ZN => maptoVGA(204));
  mapmech_t19_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t19_n_2, Q => mapmech_t19_state);
  mapmech_t19_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(204), A2 => mapmech_t19_n_1, B => n_0, C => mapmech_t19_n_0, ZN => mapmech_t19_n_2);
  mapmech_t19_g119 : ND2D0BWP7T port map(A1 => mapmech_xo7, A2 => mapmech_yo1, ZN => mapmech_t19_n_1);
  mapmech_t19_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t19_n_0);
  mapmech_t20_g68 : INVD4BWP7T port map(I => mapmech_t20_state, ZN => maptoVGA(202));
  mapmech_t20_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t20_n_2, Q => mapmech_t20_state);
  mapmech_t20_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(202), A2 => mapmech_t20_n_1, B => n_0, C => mapmech_t20_n_0, ZN => mapmech_t20_n_2);
  mapmech_t20_g119 : ND2D0BWP7T port map(A1 => mapmech_xo8, A2 => mapmech_yo1, ZN => mapmech_t20_n_1);
  mapmech_t20_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t20_n_0);
  mapmech_t92_g136 : BUFFD4BWP7T port map(I => mapmech_t92_state(1), Z => maptoVGA(58));
  mapmech_t92_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t92_n_7, A2 => mapmech_t92_n_8, Z => maptoVGA(59));
  mapmech_t92_g185 : NR2XD0BWP7T port map(A1 => mapmech_t92_n_4, A2 => n_0, ZN => mapmech_t92_n_6);
  mapmech_t92_g186 : AOI21D0BWP7T port map(A1 => mapmech_t92_n_2, A2 => mapmech_t92_n_3, B => n_0, ZN => mapmech_t92_n_5);
  mapmech_t92_g187 : AOI22D0BWP7T port map(A1 => mapmech_t92_state(1), A2 => mapmech_t92_n_3, B1 => mapmech_t92_state(0), B2 => mapmech_t92_n_1, ZN => mapmech_t92_n_4);
  mapmech_t92_g188 : ND3D0BWP7T port map(A1 => mapmech_xo3, A2 => mapmech_yo8, A3 => n_105, ZN => mapmech_t92_n_3);
  mapmech_t92_g189 : ND2D1BWP7T port map(A1 => mapmech_t92_state(0), A2 => n_105, ZN => mapmech_t92_n_2);
  mapmech_t92_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t92_n_1);
  mapmech_t92_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t92_n_5, Q => mapmech_t92_state(0), QN => mapmech_t92_n_8);
  mapmech_t92_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t92_n_6, Q => mapmech_t92_state(1), QN => mapmech_t92_n_7);
  mapmech_t21_g68 : INVD4BWP7T port map(I => mapmech_t21_state, ZN => maptoVGA(200));
  mapmech_t21_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t21_n_2, Q => mapmech_t21_state);
  mapmech_t21_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(200), A2 => mapmech_t21_n_1, B => n_0, C => mapmech_t21_n_0, ZN => mapmech_t21_n_2);
  mapmech_t21_g119 : ND2D0BWP7T port map(A1 => mapmech_xo9, A2 => mapmech_yo1, ZN => mapmech_t21_n_1);
  mapmech_t21_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t21_n_0);
  mapmech_t94_g136 : BUFFD4BWP7T port map(I => mapmech_t94_state(1), Z => maptoVGA(54));
  mapmech_t94_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t94_n_7, A2 => mapmech_t94_n_8, Z => maptoVGA(55));
  mapmech_t94_g185 : NR2XD0BWP7T port map(A1 => mapmech_t94_n_4, A2 => n_0, ZN => mapmech_t94_n_6);
  mapmech_t94_g186 : AOI21D0BWP7T port map(A1 => mapmech_t94_n_2, A2 => mapmech_t94_n_3, B => n_0, ZN => mapmech_t94_n_5);
  mapmech_t94_g187 : AOI22D0BWP7T port map(A1 => mapmech_t94_state(1), A2 => mapmech_t94_n_3, B1 => mapmech_t94_state(0), B2 => mapmech_t94_n_1, ZN => mapmech_t94_n_4);
  mapmech_t94_g188 : ND3D0BWP7T port map(A1 => mapmech_xo5, A2 => mapmech_yo8, A3 => n_105, ZN => mapmech_t94_n_3);
  mapmech_t94_g189 : ND2D1BWP7T port map(A1 => mapmech_t94_state(0), A2 => n_105, ZN => mapmech_t94_n_2);
  mapmech_t94_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t94_n_1);
  mapmech_t94_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t94_n_5, Q => mapmech_t94_state(0), QN => mapmech_t94_n_8);
  mapmech_t94_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t94_n_6, Q => mapmech_t94_state(1), QN => mapmech_t94_n_7);
  mapmech_t24_g68 : INVD4BWP7T port map(I => mapmech_t24_state, ZN => maptoVGA(194));
  mapmech_t24_state_reg : DFQD1BWP7T port map(CP => clk, D => mapmech_t24_n_2, Q => mapmech_t24_state);
  mapmech_t24_g118 : AOI211XD0BWP7T port map(A1 => maptoVGA(194), A2 => mapmech_t24_n_1, B => n_0, C => mapmech_t24_n_0, ZN => mapmech_t24_n_2);
  mapmech_t24_g119 : ND2D0BWP7T port map(A1 => mapmech_xo1, A2 => mapmech_yo2, ZN => mapmech_t24_n_1);
  mapmech_t24_g120 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t24_n_0);
  mapmech_t96_g136 : BUFFD4BWP7T port map(I => mapmech_t96_state(1), Z => maptoVGA(50));
  mapmech_t96_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t96_n_7, A2 => mapmech_t96_n_9, Z => maptoVGA(51));
  mapmech_t96_g185 : NR2XD0BWP7T port map(A1 => mapmech_t96_n_4, A2 => n_0, ZN => mapmech_t96_n_6);
  mapmech_t96_g186 : AOI21D0BWP7T port map(A1 => mapmech_t96_n_2, A2 => mapmech_t96_n_3, B => n_0, ZN => mapmech_t96_n_5);
  mapmech_t96_g187 : AOI22D0BWP7T port map(A1 => mapmech_t96_state(1), A2 => mapmech_t96_n_3, B1 => mapmech_t96_state(0), B2 => mapmech_t96_n_1, ZN => mapmech_t96_n_4);
  mapmech_t96_g188 : ND3D0BWP7T port map(A1 => mapmech_xo7, A2 => mapmech_yo8, A3 => n_105, ZN => mapmech_t96_n_3);
  mapmech_t96_g189 : ND2D1BWP7T port map(A1 => mapmech_t96_state(0), A2 => n_105, ZN => mapmech_t96_n_2);
  mapmech_t96_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t96_n_1);
  mapmech_t96_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t96_n_5, Q => mapmech_t96_state(0), QN => mapmech_t96_n_9);
  mapmech_t96_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t96_n_6, Q => mapmech_t96_state(1), QN => mapmech_t96_n_7);
  mapmech_t26_g136 : BUFFD4BWP7T port map(I => mapmech_t26_state(1), Z => maptoVGA(190));
  mapmech_t26_g141 : CKAN2D8BWP7T port map(A1 => mapmech_t26_n_7, A2 => mapmech_t26_n_8, Z => maptoVGA(191));
  mapmech_t26_g185 : NR2XD0BWP7T port map(A1 => mapmech_t26_n_4, A2 => n_0, ZN => mapmech_t26_n_6);
  mapmech_t26_g186 : AOI21D0BWP7T port map(A1 => mapmech_t26_n_2, A2 => mapmech_t26_n_3, B => n_0, ZN => mapmech_t26_n_5);
  mapmech_t26_g187 : AOI22D0BWP7T port map(A1 => mapmech_t26_state(1), A2 => mapmech_t26_n_3, B1 => mapmech_t26_state(0), B2 => mapmech_t26_n_1, ZN => mapmech_t26_n_4);
  mapmech_t26_g188 : ND3D0BWP7T port map(A1 => mapmech_xo3, A2 => mapmech_yo2, A3 => n_105, ZN => mapmech_t26_n_3);
  mapmech_t26_g189 : ND2D1BWP7T port map(A1 => mapmech_t26_state(0), A2 => n_105, ZN => mapmech_t26_n_2);
  mapmech_t26_drc_bufs192 : INVD0BWP7T port map(I => n_105, ZN => mapmech_t26_n_1);
  mapmech_t26_state_reg_0 : DFD1BWP7T port map(CP => clk, D => mapmech_t26_n_5, Q => mapmech_t26_state(0), QN => mapmech_t26_n_8);
  mapmech_t26_state_reg_1 : DFD1BWP7T port map(CP => clk, D => mapmech_t26_n_6, Q => mapmech_t26_state(1), QN => mapmech_t26_n_7);
  tie_0_cell : TIELBWP7T port map(ZN => maptoVGA(217));
  tie_1_cell : TIEHBWP7T port map(Z => maptoVGA(241));

end synthesised;
