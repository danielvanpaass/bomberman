library IEEE;
use IEEE.std_logic_1164.ALL;

entity last_bomb_tb is
end last_bomb_tb;

