library IEEE;
use IEEE.std_logic_1164.ALL;

entity obstacle_map_tb is
end obstacle_map_tb;

