configuration vga_controller_behaviour_cfg of vga_controller is
   for behaviour
   end for;
end vga_controller_behaviour_cfg;
