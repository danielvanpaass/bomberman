configuration sprites_tb_behaviour_cfg of sprites_tb is
   for behaviour
      for all: sprites use configuration work.sprites_behaviour_cfg;
      end for;
   end for;
end sprites_tb_behaviour_cfg;
