library IEEE;
use IEEE.std_logic_1164.ALL;

entity sprites_tb is
end sprites_tb;

