library IEEE;
use IEEE.std_logic_1164.ALL;

entity tile_stdempty_tb is
end tile_stdempty_tb;

