library IEEE;
use IEEE.std_logic_1164.ALL;

entity test_tb is
end test_tb;

