library IEEE;
use IEEE.std_logic_1164.ALL;

entity toplvl_coor_tb is
end toplvl_coor_tb;

