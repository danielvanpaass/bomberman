configuration hitbox_synthesised_cfg of hitbox is
   for synthesised
   end for;
end hitbox_synthesised_cfg;
