library IEEE;
use IEEE.std_logic_1164.ALL;

entity buff_tb is
end buff_tb;

