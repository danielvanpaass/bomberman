configuration hitbox_hitbox_behaviour_cfg of hitbox is
   for hitbox_behaviour
   end for;
end hitbox_hitbox_behaviour_cfg;
