configuration buff_behaviour_cfg of buff is
   for behaviour
      for all: reg use configuration work.reg_behaviour_cfg;
      end for;
   end for;
end buff_behaviour_cfg;
