library IEEE;
use IEEE.std_logic_1164.ALL;

entity bombhandling_tb is
end bombhandling_tb;

