LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
ARCHITECTURE behaviour OF hitbox_tb IS
 COMPONENT hitbox
  PORT (
   clk              : IN std_logic;
   reset            : IN std_logic;
   walls_and_crates : IN std_logic_vector(120 DOWNTO 0);
   bomb_x_a         : IN std_logic_vector(3 DOWNTO 0);
   bomb_y_a         : IN std_logic_vector(3 DOWNTO 0);
   bomb_x_b         : IN std_logic_vector(3 DOWNTO 0);
   bomb_y_b         : IN std_logic_vector(3 DOWNTO 0);
   bomb_x_c         : IN std_logic_vector(3 DOWNTO 0);
   bomb_y_c         : IN std_logic_vector(3 DOWNTO 0);
   bomb_x_d         : IN std_logic_vector(3 DOWNTO 0);
   bomb_y_d         : IN std_logic_vector(3 DOWNTO 0);
   bomb_x_e         : IN std_logic_vector(3 DOWNTO 0);
   bomb_y_e         : IN std_logic_vector(3 DOWNTO 0);
   bomb_x_f         : IN std_logic_vector(3 DOWNTO 0);
   bomb_y_f         : IN std_logic_vector(3 DOWNTO 0);
   bomb_x_g         : IN std_logic_vector(3 DOWNTO 0);
   bomb_y_g         : IN std_logic_vector(3 DOWNTO 0);
   bomb_x_h         : IN std_logic_vector(3 DOWNTO 0);
   bomb_y_h         : IN std_logic_vector(3 DOWNTO 0);
   bomb_a_active    : IN std_logic;
   bomb_b_active    : IN std_logic;
   bomb_c_active    : IN std_logic;
   bomb_d_active    : IN std_logic;
   bomb_e_active    : IN std_logic;
   bomb_f_active    : IN std_logic;
   bomb_g_active    : IN std_logic;
   bomb_h_active    : IN std_logic;
   up_p1            : IN std_logic;
   right_p1         : IN std_logic;
   down_p1          : IN std_logic;
   left_p1          : IN std_logic;
   up_p2            : IN std_logic;
   right_p2         : IN std_logic;
   down_p2          : IN std_logic;
   left_p2          : IN std_logic;
   x_p1             : OUT std_logic_vector(3 DOWNTO 0);
   y_p1             : OUT std_logic_vector(3 DOWNTO 0);
   x_p2             : OUT std_logic_vector(3 DOWNTO 0);
   y_p2             : OUT std_logic_vector(3 DOWNTO 0)
  );
 END COMPONENT;
 SIGNAL clk              : std_logic;
 SIGNAL reset            : std_logic;
 SIGNAL walls_and_crates : std_logic_vector(120 DOWNTO 0);
 SIGNAL bomb_x_a         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_y_a         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_x_b         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_y_b         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_x_c         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_y_c         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_x_d         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_y_d         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_x_e         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_y_e         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_x_f         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_y_f         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_x_g         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_y_g         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_x_h         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_y_h         : std_logic_vector(3 DOWNTO 0);
 SIGNAL bomb_a_active    : std_logic;
 SIGNAL bomb_b_active    : std_logic;
 SIGNAL bomb_c_active    : std_logic;
 SIGNAL bomb_d_active    : std_logic;
 SIGNAL bomb_e_active    : std_logic;
 SIGNAL bomb_f_active    : std_logic;
 SIGNAL bomb_g_active    : std_logic;
 SIGNAL bomb_h_active    : std_logic;
 SIGNAL up_p1            : std_logic;
 SIGNAL right_p1         : std_logic;
 SIGNAL down_p1          : std_logic;
 SIGNAL left_p1          : std_logic;
 SIGNAL up_p2            : std_logic;
 SIGNAL right_p2         : std_logic;
 SIGNAL down_p2          : std_logic;
 SIGNAL left_p2          : std_logic;
 SIGNAL x_p1             : std_logic_vector(3 DOWNTO 0);
 SIGNAL y_p1             : std_logic_vector(3 DOWNTO 0);
 SIGNAL x_p2             : std_logic_vector(3 DOWNTO 0);
 SIGNAL y_p2             : std_logic_vector(3 DOWNTO 0);
BEGIN
 test : hitbox
 PORT MAP(clk, reset, walls_and_crates, bomb_x_a, bomb_y_a, bomb_x_b, bomb_y_b, bomb_x_c, bomb_y_c, bomb_x_d, bomb_y_d, bomb_x_e, bomb_y_e, bomb_x_f, bomb_y_f, bomb_x_g, bomb_y_g, bomb_x_h, bomb_y_h, bomb_a_active, bomb_b_active, bomb_c_active, bomb_d_active, bomb_e_active, bomb_f_active, bomb_g_active, up_p1, right_p1, down_p1, left_p1, up_p2, right_p2, down_p2, left_p2, x_p1, y_p1, x_p2, y_p2);
 clk <= '1' AFTER 0 ns,
  '0' AFTER 0.04 ms WHEN clk /= '0' ELSE '1' AFTER 0.04 ms;
  reset <= '1' AFTER 0 ns,
   '0' AFTER 0.12 ms;
   walls_and_crates <= "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" AFTER 0 ns;
   bomb_x_a         <= "0000" AFTER 0 ns;
   bomb_y_a         <= "0000" AFTER 0 ns;
   bomb_x_b         <= "0000" AFTER 0 ns;
   bomb_y_b         <= "0000" AFTER 0 ns;
   bomb_x_c         <= "0000" AFTER 0 ns;
   bomb_y_c         <= "0000" AFTER 0 ns;
   bomb_x_d         <= "0000" AFTER 0 ns;
   bomb_y_d         <= "0000" AFTER 0 ns;
   bomb_x_e         <= "0000" AFTER 0 ns;
   bomb_y_e         <= "0000" AFTER 0 ns;
   bomb_x_f         <= "0000" AFTER 0 ns;
   bomb_y_f         <= "0000" AFTER 0 ns;
   bomb_x_g         <= "0000" AFTER 0 ns;
   bomb_y_g         <= "0000" AFTER 0 ns;
   bomb_x_h         <= "0000" AFTER 0 ns;
   bomb_y_h         <= "0000" AFTER 0 ns;
   bomb_a_active    <= '0' AFTER 0 ns;
   bomb_b_active    <= '0' AFTER 0 ns;
   bomb_c_active    <= '0' AFTER 0 ns;
   bomb_d_active    <= '0' AFTER 0 ns;
   bomb_e_active    <= '0' AFTER 0 ns;
   bomb_f_active    <= '0' AFTER 0 ns;
   bomb_g_active    <= '0' AFTER 0 ns;
   bomb_h_active    <= '0' AFTER 0 ns;
   up_p1            <= '0' AFTER 0 ns;
   right_p1         <= '0' AFTER 0 ns,
    '1' AFTER 4 ms;
    down_p1  <= '0' AFTER 0 ns;
    left_p1  <= '0' AFTER 0 ns;
    up_p2    <= '0' AFTER 0 ns;
    right_p2 <= '0' AFTER 0 ns;
    down_p2  <= '0' AFTER 0 ns;
    left_p2  <= '0' AFTER 0 ns,
     '1' AFTER 3 ms;
END behaviour;
