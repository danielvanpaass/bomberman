configuration tile_stdempty_tb_behaviour_cfg of tile_stdempty_tb is
   for behaviour
      for all: tile_stdempty use configuration work.tile_stdempty_behaviour_cfg;
      end for;
   end for;
end tile_stdempty_tb_behaviour_cfg;
