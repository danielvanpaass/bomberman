configuration uneven_bits_tb_behaviour_cfg of uneven_bits_tb is
   for behaviour
      for all: uneven_bits use configuration work.uneven_bits_behaviour_cfg;
      end for;
   end for;
end uneven_bits_tb_behaviour_cfg;
