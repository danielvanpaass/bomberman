configuration obstacle_map_behaviour_cfg of obstacle_map is
   for behaviour
      for all: uneven_bits use configuration work.uneven_bits_behaviour_cfg;
      end for;
   end for;
end obstacle_map_behaviour_cfg;
