library IEEE;
use IEEE.std_logic_1164.ALL;

entity selector_tb is
end selector_tb;

