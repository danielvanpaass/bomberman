library IEEE;
use IEEE.std_logic_1164.ALL;

entity sprites is
   port(clk : in std_logic;
reset : in std_logic;
victory : in std_logic;
playground_y0 : in  std_logic_vector(21 downto 0);
playground_y1 : in  std_logic_vector(21 downto 0);
playground_y2 : in  std_logic_vector(21 downto 0);
playground_y3 : in  std_logic_vector(21 downto 0);
playground_y4 : in  std_logic_vector(21 downto 0);
playground_y5 : in  std_logic_vector(21 downto 0);
playground_y6 : in  std_logic_vector(21 downto 0);
playground_y7 : in  std_logic_vector(21 downto 0);
playground_y8 : in  std_logic_vector(21 downto 0);
playground_y9 : in  std_logic_vector(21 downto 0);
playground_y10 : in  std_logic_vector(21 downto 0);
        x_p1          : in  std_logic_vector(3 downto 0);
        y_p1          : in  std_logic_vector(3 downto 0);
       x_p2          : in  std_logic_vector(3 downto 0);
       y_p2          : in  std_logic_vector(3 downto 0);
        x_bomb_a      : in  std_logic_vector(3 downto 0);
        y_bomb_a      : in  std_logic_vector(3 downto 0);
        bomb_a_enable : in  std_logic;
        x_bomb_b      : in  std_logic_vector(3 downto 0);
        y_bomb_b      : in  std_logic_vector(3 downto 0);
        bomb_b_enable : in  std_logic;
        x_bomb_c      : in  std_logic_vector(3 downto 0);
        y_bomb_c      : in  std_logic_vector(3 downto 0);
        bomb_c_enable : in  std_logic;
        x_bomb_d      : in  std_logic_vector(3 downto 0);
        y_bomb_d      : in  std_logic_vector(3 downto 0);
        bomb_d_enable : in  std_logic;
        x_bomb_e      : in  std_logic_vector(3 downto 0);
        y_bomb_e      : in  std_logic_vector(3 downto 0);
        bomb_e_enable : in  std_logic;
        x_bomb_f      : in  std_logic_vector(3 downto 0);
        y_bomb_f      : in  std_logic_vector(3 downto 0);
        bomb_f_enable : in  std_logic;
        x_bomb_g      : in  std_logic_vector(3 downto 0);
        y_bomb_g      : in  std_logic_vector(3 downto 0);
        bomb_g_enable : in  std_logic;
        x_bomb_h      : in  std_logic_vector(3 downto 0);
        y_bomb_h      : in  std_logic_vector(3 downto 0);
        bomb_h_enable : in  std_logic;
        x_map         : in  std_logic_vector(3 downto 0);
        y_map         : in  std_logic_vector(3 downto 0);
        input_h_map         : in  std_logic_vector(4 downto 0);
        input_v_map         : in  std_logic_vector(5 downto 0);
        rgb           : out std_logic_vector(2 downto 0));
end sprites;

