
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of playground is

  component INVD1BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component INVD4BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component DFQD1BWP7T
    port(CP, D : in std_logic; Q : out std_logic);
  end component;

  component AOI211XD0BWP7T
    port(A1, A2, B, C : in std_logic; ZN : out std_logic);
  end component;

  component ND2D0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component INVD0BWP7T
    port(I : in std_logic; ZN : out std_logic);
  end component;

  component BUFFD4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;

  component AN2D4BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component NR2XD0BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component AOI21D0BWP7T
    port(A1, A2, B : in std_logic; ZN : out std_logic);
  end component;

  component AOI22D0BWP7T
    port(A1, A2, B1, B2 : in std_logic; ZN : out std_logic);
  end component;

  component ND3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component ND2D1BWP7T
    port(A1, A2 : in std_logic; ZN : out std_logic);
  end component;

  component DFD1BWP7T
    port(CP, D : in std_logic; Q, QN : out std_logic);
  end component;

  component INR2XD0BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component NR3D0BWP7T
    port(A1, A2, A3 : in std_logic; ZN : out std_logic);
  end component;

  component IND2D1BWP7T
    port(A1, B1 : in std_logic; ZN : out std_logic);
  end component;

  component OR2D1BWP7T
    port(A1, A2 : in std_logic; Z : out std_logic);
  end component;

  component TIELBWP7T
    port(ZN : out std_logic);
  end component;

  component TIEHBWP7T
    port(Z : out std_logic);
  end component;

  signal t63_state : std_logic_vector(1 downto 0);
  signal t64_state : std_logic_vector(1 downto 0);
  signal t65_state : std_logic_vector(1 downto 0);
  signal t68_state : std_logic_vector(1 downto 0);
  signal t70_state : std_logic_vector(1 downto 0);
  signal t74_state : std_logic_vector(1 downto 0);
  signal t76_state : std_logic_vector(1 downto 0);
  signal t80_state : std_logic_vector(1 downto 0);
  signal t81_state : std_logic_vector(1 downto 0);
  signal t82_state : std_logic_vector(1 downto 0);
  signal t83_state : std_logic_vector(1 downto 0);
  signal t84_state : std_logic_vector(1 downto 0);
  signal t104_state : std_logic_vector(1 downto 0);
  signal t85_state : std_logic_vector(1 downto 0);
  signal t105_state : std_logic_vector(1 downto 0);
  signal t86_state : std_logic_vector(1 downto 0);
  signal t106_state : std_logic_vector(1 downto 0);
  signal t92_state : std_logic_vector(1 downto 0);
  signal t94_state : std_logic_vector(1 downto 0);
  signal t96_state : std_logic_vector(1 downto 0);
  signal t26_state : std_logic_vector(1 downto 0);
  signal t28_state : std_logic_vector(1 downto 0);
  signal t30_state : std_logic_vector(1 downto 0);
  signal t36_state : std_logic_vector(1 downto 0);
  signal t37_state : std_logic_vector(1 downto 0);
  signal t38_state : std_logic_vector(1 downto 0);
  signal t39_state : std_logic_vector(1 downto 0);
  signal t40_state : std_logic_vector(1 downto 0);
  signal t41_state : std_logic_vector(1 downto 0);
  signal t42_state : std_logic_vector(1 downto 0);
  signal t46_state : std_logic_vector(1 downto 0);
  signal t48_state : std_logic_vector(1 downto 0);
  signal t52_state : std_logic_vector(1 downto 0);
  signal t54_state : std_logic_vector(1 downto 0);
  signal t57_state : std_logic_vector(1 downto 0);
  signal t58_state : std_logic_vector(1 downto 0);
  signal t59_state : std_logic_vector(1 downto 0);
  signal n_126, n_128, n_141, n_142, t13_n_1 : std_logic;
  signal t13_n_2, t13_n_3, t13_state, t14_n_1, t14_n_2 : std_logic;
  signal t14_n_3, t14_state, t15_n_1, t15_n_2, t15_n_3 : std_logic;
  signal t15_state, t19_n_1, t19_n_2, t19_n_3, t19_state : std_logic;
  signal t20_n_1, t20_n_2, t20_n_3, t20_state, t21_n_1 : std_logic;
  signal t21_n_2, t21_n_3, t21_state, t24_n_1, t24_n_2 : std_logic;
  signal t24_n_3, t24_state, t26_n_2, t26_n_3, t26_n_4 : std_logic;
  signal t26_n_5, t26_n_6, t26_n_7, t26_n_8, t26_n_9 : std_logic;
  signal t26_n_10, t28_n_2, t28_n_3, t28_n_4, t28_n_5 : std_logic;
  signal t28_n_6, t28_n_7, t28_n_8, t28_n_9, t28_n_10 : std_logic;
  signal t30_n_3, t30_n_4, t30_n_5, t30_n_6, t30_n_7 : std_logic;
  signal t30_n_8, t30_n_9, t30_n_10, t32_n_1, t32_n_2 : std_logic;
  signal t32_n_3, t32_state, t35_n_1, t35_n_2, t35_n_3 : std_logic;
  signal t35_state, t36_n_2, t36_n_3, t36_n_4, t36_n_5 : std_logic;
  signal t36_n_6, t36_n_7, t36_n_8, t36_n_9, t36_n_10 : std_logic;
  signal t37_n_3, t37_n_4, t37_n_5, t37_n_6, t37_n_7 : std_logic;
  signal t37_n_8, t37_n_9, t37_n_10, t38_n_2, t38_n_3 : std_logic;
  signal t38_n_4, t38_n_5, t38_n_6, t38_n_7, t38_n_8 : std_logic;
  signal t38_n_9, t38_n_10, t39_n_0, t39_n_1, t39_n_2 : std_logic;
  signal t39_n_3, t39_n_4, t39_n_5, t39_n_6, t39_n_7 : std_logic;
  signal t39_n_8, t39_n_9, t39_n_10, t40_n_2, t40_n_3 : std_logic;
  signal t40_n_4, t40_n_5, t40_n_6, t40_n_7, t40_n_8 : std_logic;
  signal t40_n_9, t40_n_10, t41_n_3, t41_n_4, t41_n_5 : std_logic;
  signal t41_n_6, t41_n_7, t41_n_8, t41_n_9, t41_n_10 : std_logic;
  signal t42_n_0, t42_n_1, t42_n_2, t42_n_3, t42_n_4 : std_logic;
  signal t42_n_5, t42_n_6, t42_n_7, t42_n_8, t42_n_9 : std_logic;
  signal t42_n_10, t43_n_1, t43_n_2, t43_n_3, t43_state : std_logic;
  signal t46_n_2, t46_n_3, t46_n_4, t46_n_5, t46_n_6 : std_logic;
  signal t46_n_7, t46_n_8, t46_n_9, t46_n_11, t48_n_3 : std_logic;
  signal t48_n_4, t48_n_5, t48_n_6, t48_n_7, t48_n_8 : std_logic;
  signal t48_n_9, t48_n_10, t50_n_1, t50_n_2, t50_n_3 : std_logic;
  signal t50_state, t52_n_0, t52_n_1, t52_n_2, t52_n_3 : std_logic;
  signal t52_n_4, t52_n_5, t52_n_6, t52_n_7, t52_n_8 : std_logic;
  signal t52_n_9, t52_n_11, t54_n_2, t54_n_3, t54_n_4 : std_logic;
  signal t54_n_5, t54_n_6, t54_n_7, t54_n_8, t54_n_9 : std_logic;
  signal t54_n_11, t57_n_3, t57_n_4, t57_n_5, t57_n_6 : std_logic;
  signal t57_n_7, t57_n_8, t57_n_9, t57_n_11, t58_n_0 : std_logic;
  signal t58_n_1, t58_n_2, t58_n_3, t58_n_4, t58_n_5 : std_logic;
  signal t58_n_6, t58_n_7, t58_n_8, t58_n_9, t58_n_10 : std_logic;
  signal t59_n_2, t59_n_3, t59_n_4, t59_n_5, t59_n_6 : std_logic;
  signal t59_n_7, t59_n_8, t59_n_9, t59_n_11, t60_n_1 : std_logic;
  signal t60_n_2, t60_n_3, t60_state, t61_n_1, t61_n_2 : std_logic;
  signal t61_n_3, t61_state, t62_n_1, t62_n_2, t62_n_3 : std_logic;
  signal t62_state, t63_n_2, t63_n_3, t63_n_4, t63_n_5 : std_logic;
  signal t63_n_6, t63_n_7, t63_n_8, t63_n_9, t63_n_10 : std_logic;
  signal t64_n_2, t64_n_3, t64_n_4, t64_n_5, t64_n_6 : std_logic;
  signal t64_n_7, t64_n_8, t64_n_9, t64_n_10, t65_n_3 : std_logic;
  signal t65_n_4, t65_n_5, t65_n_6, t65_n_7, t65_n_8 : std_logic;
  signal t65_n_9, t65_n_11, t68_n_3, t68_n_4, t68_n_5 : std_logic;
  signal t68_n_6, t68_n_7, t68_n_8, t68_n_9, t68_n_10 : std_logic;
  signal t70_n_0, t70_n_1, t70_n_2, t70_n_3, t70_n_4 : std_logic;
  signal t70_n_5, t70_n_6, t70_n_7, t70_n_8, t70_n_9 : std_logic;
  signal t70_n_10, t72_n_1, t72_n_2, t72_n_3, t72_state : std_logic;
  signal t74_n_0, t74_n_1, t74_n_3, t74_n_4, t74_n_5 : std_logic;
  signal t74_n_6, t74_n_7, t74_n_8, t74_n_9, t74_n_10 : std_logic;
  signal t76_n_2, t76_n_3, t76_n_4, t76_n_5, t76_n_6 : std_logic;
  signal t76_n_7, t76_n_8, t76_n_9, t76_n_10, t79_n_1 : std_logic;
  signal t79_n_2, t79_n_3, t79_state, t80_n_2, t80_n_3 : std_logic;
  signal t80_n_4, t80_n_5, t80_n_6, t80_n_7, t80_n_8 : std_logic;
  signal t80_n_9, t80_n_10, t81_n_0, t81_n_1, t81_n_3 : std_logic;
  signal t81_n_4, t81_n_5, t81_n_6, t81_n_7, t81_n_8 : std_logic;
  signal t81_n_9, t81_n_10, t82_n_2, t82_n_3, t82_n_4 : std_logic;
  signal t82_n_5, t82_n_6, t82_n_7, t82_n_8, t82_n_9 : std_logic;
  signal t82_n_10, t83_n_2, t83_n_3, t83_n_4, t83_n_5 : std_logic;
  signal t83_n_6, t83_n_7, t83_n_8, t83_n_9, t83_n_11 : std_logic;
  signal t84_n_0, t84_n_1, t84_n_2, t84_n_3, t84_n_4 : std_logic;
  signal t84_n_5, t84_n_6, t84_n_7, t84_n_8, t84_n_9 : std_logic;
  signal t84_n_10, t85_n_0, t85_n_1, t85_n_3, t85_n_4 : std_logic;
  signal t85_n_5, t85_n_6, t85_n_7, t85_n_8, t85_n_9 : std_logic;
  signal t85_n_10, t86_n_2, t86_n_3, t86_n_4, t86_n_5 : std_logic;
  signal t86_n_6, t86_n_7, t86_n_8, t86_n_9, t86_n_10 : std_logic;
  signal t87_n_1, t87_n_2, t87_n_3, t87_state, t90_n_1 : std_logic;
  signal t90_n_2, t90_n_3, t90_state, t92_n_3, t92_n_4 : std_logic;
  signal t92_n_5, t92_n_6, t92_n_7, t92_n_8, t92_n_9 : std_logic;
  signal t92_n_11, t94_n_2, t94_n_3, t94_n_4, t94_n_5 : std_logic;
  signal t94_n_6, t94_n_7, t94_n_8, t94_n_9, t94_n_10 : std_logic;
  signal t96_n_2, t96_n_3, t96_n_4, t96_n_5, t96_n_6 : std_logic;
  signal t96_n_7, t96_n_8, t96_n_9, t96_n_11, t98_n_1 : std_logic;
  signal t98_n_2, t98_n_3, t98_state, t101_n_1, t101_n_2 : std_logic;
  signal t101_n_3, t101_state, t102_n_1, t102_n_2, t102_n_3 : std_logic;
  signal t102_state, t103_n_1, t103_n_2, t103_n_3, t103_state : std_logic;
  signal t104_n_2, t104_n_3, t104_n_4, t104_n_5, t104_n_6 : std_logic;
  signal t104_n_7, t104_n_8, t104_n_9, t104_n_11, t105_n_3 : std_logic;
  signal t105_n_4, t105_n_5, t105_n_6, t105_n_7, t105_n_8 : std_logic;
  signal t105_n_9, t105_n_11, t106_n_0, t106_n_1, t106_n_2 : std_logic;
  signal t106_n_3, t106_n_4, t106_n_5, t106_n_6, t106_n_7 : std_logic;
  signal t106_n_8, t106_n_9, t106_n_10, t107_n_1, t107_n_2 : std_logic;
  signal t107_n_3, t107_state, t108_n_1, t108_n_2, t108_n_3 : std_logic;
  signal t108_state, t109_n_1, t109_n_2, t109_n_3, t109_state : std_logic;
  signal tt16_n_1, tt16_n_2, tt16_n_3, tt16_state, tt17_n_1 : std_logic;
  signal tt17_n_2, tt17_n_3, tt17_state, tt18_n_1, tt18_n_2 : std_logic;
  signal tt18_n_3, tt18_state, xo1, xo2, xo3 : std_logic;
  signal xo4, xo5, xo6, xo7, xo8 : std_logic;
  signal xo9, xyconv_n_1, xyconv_n_2, xyconv_n_3, xyconv_n_4 : std_logic;
  signal xyconv_n_5, xyconv_n_6, xyconv_n_7, xyconv_n_8, xyconv_n_10 : std_logic;
  signal xyconv_n_11, xyconv_n_12, xyconv_n_14, xyconv_n_15, xyconv_n_16 : std_logic;
  signal yo1, yo2, yo3, yo4, yo5 : std_logic;
  signal yo6, yo7, yo8, yo9 : std_logic;

begin

  y10(0) <= y0(21);
  y10(1) <= y0(21);
  y10(2) <= y0(21);
  y10(3) <= y0(21);
  y10(4) <= y0(21);
  y10(5) <= y0(21);
  y10(6) <= y0(21);
  y10(7) <= y0(21);
  y10(8) <= y0(21);
  y10(9) <= y0(21);
  y10(10) <= y0(21);
  y10(11) <= y0(21);
  y10(12) <= y0(21);
  y10(13) <= y0(21);
  y10(14) <= y0(21);
  y10(15) <= y0(21);
  y10(16) <= y0(21);
  y10(17) <= y0(21);
  y10(18) <= y0(21);
  y10(19) <= y0(21);
  y10(20) <= y0(21);
  y10(21) <= y0(21);
  y9(0) <= y0(21);
  y9(1) <= y0(21);
  y9(3) <= y1(19);
  y9(5) <= y1(19);
  y9(7) <= y1(19);
  y9(15) <= y1(19);
  y9(17) <= y1(19);
  y9(19) <= y1(19);
  y9(20) <= y0(21);
  y9(21) <= y0(21);
  y8(0) <= y0(21);
  y8(1) <= y0(21);
  y8(3) <= y1(19);
  y8(4) <= y0(21);
  y8(5) <= y0(21);
  y8(8) <= y0(21);
  y8(9) <= y0(21);
  y8(12) <= y0(21);
  y8(13) <= y0(21);
  y8(16) <= y0(21);
  y8(17) <= y0(21);
  y8(19) <= y1(19);
  y8(20) <= y0(21);
  y8(21) <= y0(21);
  y7(0) <= y0(21);
  y7(1) <= y0(21);
  y7(3) <= y1(19);
  y7(19) <= y1(19);
  y7(20) <= y0(21);
  y7(21) <= y0(21);
  y6(0) <= y0(21);
  y6(1) <= y0(21);
  y6(4) <= y0(21);
  y6(5) <= y0(21);
  y6(8) <= y0(21);
  y6(9) <= y0(21);
  y6(11) <= y1(19);
  y6(12) <= y0(21);
  y6(13) <= y0(21);
  y6(16) <= y0(21);
  y6(17) <= y0(21);
  y6(20) <= y0(21);
  y6(21) <= y0(21);
  y5(0) <= y0(21);
  y5(1) <= y0(21);
  y5(9) <= y1(19);
  y5(11) <= y1(19);
  y5(13) <= y1(19);
  y5(20) <= y0(21);
  y5(21) <= y0(21);
  y4(0) <= y0(21);
  y4(1) <= y0(21);
  y4(4) <= y0(21);
  y4(5) <= y0(21);
  y4(8) <= y0(21);
  y4(9) <= y0(21);
  y4(11) <= y1(19);
  y4(12) <= y0(21);
  y4(13) <= y0(21);
  y4(16) <= y0(21);
  y4(17) <= y0(21);
  y4(20) <= y0(21);
  y4(21) <= y0(21);
  y3(0) <= y0(21);
  y3(1) <= y0(21);
  y3(3) <= y1(19);
  y3(19) <= y1(19);
  y3(20) <= y0(21);
  y3(21) <= y0(21);
  y2(0) <= y0(21);
  y2(1) <= y0(21);
  y2(3) <= y1(19);
  y2(4) <= y0(21);
  y2(5) <= y0(21);
  y2(8) <= y0(21);
  y2(9) <= y0(21);
  y2(12) <= y0(21);
  y2(13) <= y0(21);
  y2(16) <= y0(21);
  y2(17) <= y0(21);
  y2(19) <= y1(19);
  y2(20) <= y0(21);
  y2(21) <= y0(21);
  y1(0) <= y0(21);
  y1(1) <= y0(21);
  y1(3) <= y1(19);
  y1(5) <= y1(19);
  y1(7) <= y1(19);
  y1(9) <= y1(19);
  y1(11) <= y1(19);
  y1(13) <= y1(19);
  y1(15) <= y1(19);
  y1(17) <= y1(19);
  y1(20) <= y0(21);
  y1(21) <= y0(21);
  y0(0) <= y0(21);
  y0(1) <= y0(21);
  y0(2) <= y0(21);
  y0(3) <= y0(21);
  y0(4) <= y0(21);
  y0(5) <= y0(21);
  y0(6) <= y0(21);
  y0(7) <= y0(21);
  y0(8) <= y0(21);
  y0(9) <= y0(21);
  y0(10) <= y0(21);
  y0(11) <= y0(21);
  y0(12) <= y0(21);
  y0(13) <= y0(21);
  y0(14) <= y0(21);
  y0(15) <= y0(21);
  y0(16) <= y0(21);
  y0(17) <= y0(21);
  y0(18) <= y0(21);
  y0(19) <= y0(21);
  y0(20) <= y0(21);
  drc_bufs11 : INVD1BWP7T port map(I => n_128, ZN => n_126);
  drc_bufs13 : INVD1BWP7T port map(I => reset, ZN => n_128);
  drc_bufs25 : INVD1BWP7T port map(I => n_142, ZN => n_141);
  drc_bufs26 : INVD1BWP7T port map(I => lethal, ZN => n_142);
  t61_g68 : INVD4BWP7T port map(I => t61_state, ZN => y5(10));
  t61_state_reg : DFQD1BWP7T port map(CP => clk, D => t61_n_3, Q => t61_state);
  t61_g118 : AOI211XD0BWP7T port map(A1 => y5(10), A2 => t61_n_2, B => reset, C => t61_n_1, ZN => t61_n_3);
  t61_g119 : ND2D0BWP7T port map(A1 => xo5, A2 => yo5, ZN => t61_n_2);
  t61_g120 : INVD0BWP7T port map(I => n_141, ZN => t61_n_1);
  t62_g68 : INVD4BWP7T port map(I => t62_state, ZN => y5(8));
  t62_state_reg : DFQD1BWP7T port map(CP => clk, D => t62_n_3, Q => t62_state);
  t62_g118 : AOI211XD0BWP7T port map(A1 => y5(8), A2 => t62_n_2, B => n_126, C => t62_n_1, ZN => t62_n_3);
  t62_g119 : ND2D0BWP7T port map(A1 => yo5, A2 => xo6, ZN => t62_n_2);
  t62_g120 : INVD0BWP7T port map(I => lethal, ZN => t62_n_1);
  t63_g136 : BUFFD4BWP7T port map(I => t63_state(1), Z => y5(6));
  t63_g141 : AN2D4BWP7T port map(A1 => t63_n_9, A2 => t63_n_10, Z => y5(7));
  t63_g185 : NR2XD0BWP7T port map(A1 => t63_n_6, A2 => reset, ZN => t63_n_8);
  t63_g186 : AOI21D0BWP7T port map(A1 => t63_n_4, A2 => t63_n_5, B => reset, ZN => t63_n_7);
  t63_g187 : AOI22D0BWP7T port map(A1 => t63_state(1), A2 => t63_n_5, B1 => t63_state(0), B2 => t63_n_3, ZN => t63_n_6);
  t63_g188 : ND3D0BWP7T port map(A1 => xo7, A2 => yo5, A3 => t63_n_2, ZN => t63_n_5);
  t63_g189 : ND2D1BWP7T port map(A1 => t63_state(0), A2 => t63_n_2, ZN => t63_n_4);
  t63_drc_bufs : INVD0BWP7T port map(I => t63_n_3, ZN => t63_n_2);
  t63_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t63_n_3);
  t63_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t63_n_7, Q => t63_state(0), QN => t63_n_10);
  t63_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t63_n_8, Q => t63_state(1), QN => t63_n_9);
  t64_g136 : BUFFD4BWP7T port map(I => t64_state(1), Z => y5(4));
  t64_g141 : AN2D4BWP7T port map(A1 => t64_n_9, A2 => t64_n_10, Z => y5(5));
  t64_g185 : NR2XD0BWP7T port map(A1 => t64_n_6, A2 => n_126, ZN => t64_n_8);
  t64_g186 : AOI21D0BWP7T port map(A1 => t64_n_4, A2 => t64_n_5, B => n_126, ZN => t64_n_7);
  t64_g187 : AOI22D0BWP7T port map(A1 => t64_state(1), A2 => t64_n_5, B1 => t64_state(0), B2 => t64_n_3, ZN => t64_n_6);
  t64_g188 : ND3D0BWP7T port map(A1 => yo5, A2 => xo8, A3 => t64_n_2, ZN => t64_n_5);
  t64_g189 : ND2D1BWP7T port map(A1 => t64_state(0), A2 => t64_n_2, ZN => t64_n_4);
  t64_drc_bufs : INVD0BWP7T port map(I => t64_n_3, ZN => t64_n_2);
  t64_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t64_n_3);
  t64_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t64_n_7, Q => t64_state(0), QN => t64_n_10);
  t64_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t64_n_8, Q => t64_state(1), QN => t64_n_9);
  t65_g136 : BUFFD4BWP7T port map(I => t65_state(1), Z => y5(2));
  t65_g141 : AN2D4BWP7T port map(A1 => t65_n_9, A2 => t65_n_11, Z => y5(3));
  t65_g185 : NR2XD0BWP7T port map(A1 => t65_n_6, A2 => n_126, ZN => t65_n_8);
  t65_g186 : AOI21D0BWP7T port map(A1 => t65_n_4, A2 => t65_n_5, B => n_126, ZN => t65_n_7);
  t65_g187 : AOI22D0BWP7T port map(A1 => t65_state(1), A2 => t65_n_5, B1 => t65_state(0), B2 => t65_n_3, ZN => t65_n_6);
  t65_g188 : ND3D0BWP7T port map(A1 => yo5, A2 => xo9, A3 => n_141, ZN => t65_n_5);
  t65_g189 : ND2D1BWP7T port map(A1 => t65_state(0), A2 => n_141, ZN => t65_n_4);
  t65_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t65_n_3);
  t65_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t65_n_7, Q => t65_state(0), QN => t65_n_11);
  t65_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t65_n_8, Q => t65_state(1), QN => t65_n_9);
  t68_g135 : BUFFD4BWP7T port map(I => t68_state(1), Z => y6(18));
  t68_g141 : AN2D4BWP7T port map(A1 => t68_n_9, A2 => t68_n_10, Z => y6(19));
  t68_g185 : NR2XD0BWP7T port map(A1 => t68_n_6, A2 => reset, ZN => t68_n_8);
  t68_g186 : AOI21D0BWP7T port map(A1 => t68_n_4, A2 => t68_n_5, B => reset, ZN => t68_n_7);
  t68_g187 : AOI22D0BWP7T port map(A1 => t68_state(1), A2 => t68_n_5, B1 => t68_state(0), B2 => t68_n_3, ZN => t68_n_6);
  t68_g188 : ND3D0BWP7T port map(A1 => yo6, A2 => xo1, A3 => lethal, ZN => t68_n_5);
  t68_g189 : ND2D1BWP7T port map(A1 => t68_state(0), A2 => lethal, ZN => t68_n_4);
  t68_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t68_n_3);
  t68_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t68_n_7, Q => t68_state(0), QN => t68_n_10);
  t68_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t68_n_8, Q => t68_state(1), QN => t68_n_9);
  t70_g136 : BUFFD4BWP7T port map(I => t70_state(1), Z => y6(14));
  t70_g141 : AN2D4BWP7T port map(A1 => t70_n_9, A2 => t70_n_10, Z => y6(15));
  t70_g185 : NR2XD0BWP7T port map(A1 => t70_n_6, A2 => t70_n_1, ZN => t70_n_8);
  t70_g186 : AOI21D0BWP7T port map(A1 => t70_n_4, A2 => t70_n_5, B => t70_n_1, ZN => t70_n_7);
  t70_g187 : AOI22D0BWP7T port map(A1 => t70_state(1), A2 => t70_n_5, B1 => t70_state(0), B2 => t70_n_3, ZN => t70_n_6);
  t70_g188 : ND3D0BWP7T port map(A1 => xo3, A2 => yo6, A3 => t70_n_2, ZN => t70_n_5);
  t70_g189 : ND2D1BWP7T port map(A1 => t70_state(0), A2 => t70_n_2, ZN => t70_n_4);
  t70_drc_bufs : INVD0BWP7T port map(I => t70_n_3, ZN => t70_n_2);
  t70_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t70_n_3);
  t70_drc_bufs194 : INVD0BWP7T port map(I => t70_n_0, ZN => t70_n_1);
  t70_drc_bufs196 : INVD0BWP7T port map(I => reset, ZN => t70_n_0);
  t70_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t70_n_7, Q => t70_state(0), QN => t70_n_10);
  t70_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t70_n_8, Q => t70_state(1), QN => t70_n_9);
  t72_g68 : INVD4BWP7T port map(I => t72_state, ZN => y6(10));
  t72_state_reg : DFQD1BWP7T port map(CP => clk, D => t72_n_3, Q => t72_state);
  t72_g118 : AOI211XD0BWP7T port map(A1 => y6(10), A2 => t72_n_2, B => n_126, C => t72_n_1, ZN => t72_n_3);
  t72_g119 : ND2D0BWP7T port map(A1 => xo5, A2 => yo6, ZN => t72_n_2);
  t72_g120 : INVD0BWP7T port map(I => lethal, ZN => t72_n_1);
  t74_g135 : BUFFD4BWP7T port map(I => t74_state(1), Z => y6(6));
  t74_g141 : AN2D4BWP7T port map(A1 => t74_n_9, A2 => t74_n_10, Z => y6(7));
  t74_g185 : NR2XD0BWP7T port map(A1 => t74_n_6, A2 => t74_n_1, ZN => t74_n_8);
  t74_g186 : AOI21D0BWP7T port map(A1 => t74_n_4, A2 => t74_n_5, B => t74_n_1, ZN => t74_n_7);
  t74_g187 : AOI22D0BWP7T port map(A1 => t74_state(1), A2 => t74_n_5, B1 => t74_state(0), B2 => t74_n_3, ZN => t74_n_6);
  t74_g188 : ND3D0BWP7T port map(A1 => xo7, A2 => yo6, A3 => n_141, ZN => t74_n_5);
  t74_g189 : ND2D1BWP7T port map(A1 => t74_state(0), A2 => n_141, ZN => t74_n_4);
  t74_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t74_n_3);
  t74_drc_bufs194 : INVD0BWP7T port map(I => t74_n_0, ZN => t74_n_1);
  t74_drc_bufs196 : INVD0BWP7T port map(I => reset, ZN => t74_n_0);
  t74_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t74_n_7, Q => t74_state(0), QN => t74_n_10);
  t74_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t74_n_8, Q => t74_state(1), QN => t74_n_9);
  t76_g135 : BUFFD4BWP7T port map(I => t76_state(1), Z => y6(2));
  t76_g141 : AN2D4BWP7T port map(A1 => t76_n_9, A2 => t76_n_10, Z => y6(3));
  t76_g185 : NR2XD0BWP7T port map(A1 => t76_n_6, A2 => n_126, ZN => t76_n_8);
  t76_g186 : AOI21D0BWP7T port map(A1 => t76_n_4, A2 => t76_n_5, B => n_126, ZN => t76_n_7);
  t76_g187 : AOI22D0BWP7T port map(A1 => t76_state(1), A2 => t76_n_5, B1 => t76_state(0), B2 => t76_n_3, ZN => t76_n_6);
  t76_g188 : ND3D0BWP7T port map(A1 => yo6, A2 => xo9, A3 => t76_n_2, ZN => t76_n_5);
  t76_g189 : ND2D1BWP7T port map(A1 => t76_state(0), A2 => t76_n_2, ZN => t76_n_4);
  t76_drc_bufs : INVD0BWP7T port map(I => t76_n_3, ZN => t76_n_2);
  t76_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t76_n_3);
  t76_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t76_n_7, Q => t76_state(0), QN => t76_n_10);
  t76_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t76_n_8, Q => t76_state(1), QN => t76_n_9);
  t79_g68 : INVD4BWP7T port map(I => t79_state, ZN => y7(18));
  t79_state_reg : DFQD1BWP7T port map(CP => clk, D => t79_n_3, Q => t79_state);
  t79_g118 : AOI211XD0BWP7T port map(A1 => y7(18), A2 => t79_n_2, B => reset, C => t79_n_1, ZN => t79_n_3);
  t79_g119 : ND2D0BWP7T port map(A1 => yo7, A2 => xo1, ZN => t79_n_2);
  t79_g120 : INVD0BWP7T port map(I => lethal, ZN => t79_n_1);
  t80_g136 : BUFFD4BWP7T port map(I => t80_state(1), Z => y7(16));
  t80_g141 : AN2D4BWP7T port map(A1 => t80_n_9, A2 => t80_n_10, Z => y7(17));
  t80_g185 : NR2XD0BWP7T port map(A1 => t80_n_6, A2 => n_126, ZN => t80_n_8);
  t80_g186 : AOI21D0BWP7T port map(A1 => t80_n_4, A2 => t80_n_5, B => n_126, ZN => t80_n_7);
  t80_g187 : AOI22D0BWP7T port map(A1 => t80_state(1), A2 => t80_n_5, B1 => t80_state(0), B2 => t80_n_3, ZN => t80_n_6);
  t80_g188 : ND3D0BWP7T port map(A1 => yo7, A2 => xo2, A3 => t80_n_2, ZN => t80_n_5);
  t80_g189 : ND2D1BWP7T port map(A1 => t80_state(0), A2 => t80_n_2, ZN => t80_n_4);
  t80_drc_bufs : INVD0BWP7T port map(I => t80_n_3, ZN => t80_n_2);
  t80_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t80_n_3);
  t80_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t80_n_7, Q => t80_state(0), QN => t80_n_10);
  t80_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t80_n_8, Q => t80_state(1), QN => t80_n_9);
  t81_g136 : BUFFD4BWP7T port map(I => t81_state(1), Z => y7(14));
  t81_g141 : AN2D4BWP7T port map(A1 => t81_n_9, A2 => t81_n_10, Z => y7(15));
  t81_g185 : NR2XD0BWP7T port map(A1 => t81_n_6, A2 => t81_n_1, ZN => t81_n_8);
  t81_g186 : AOI21D0BWP7T port map(A1 => t81_n_4, A2 => t81_n_5, B => t81_n_1, ZN => t81_n_7);
  t81_g187 : AOI22D0BWP7T port map(A1 => t81_state(1), A2 => t81_n_5, B1 => t81_state(0), B2 => t81_n_3, ZN => t81_n_6);
  t81_g188 : ND3D0BWP7T port map(A1 => yo7, A2 => xo3, A3 => n_141, ZN => t81_n_5);
  t81_g189 : ND2D1BWP7T port map(A1 => t81_state(0), A2 => n_141, ZN => t81_n_4);
  t81_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t81_n_3);
  t81_drc_bufs194 : INVD0BWP7T port map(I => t81_n_0, ZN => t81_n_1);
  t81_drc_bufs196 : INVD0BWP7T port map(I => reset, ZN => t81_n_0);
  t81_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t81_n_7, Q => t81_state(0), QN => t81_n_10);
  t81_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t81_n_8, Q => t81_state(1), QN => t81_n_9);
  t101_g68 : INVD4BWP7T port map(I => t101_state, ZN => y9(18));
  t101_state_reg : DFQD1BWP7T port map(CP => clk, D => t101_n_3, Q => t101_state);
  t101_g118 : AOI211XD0BWP7T port map(A1 => y9(18), A2 => t101_n_2, B => n_126, C => t101_n_1, ZN => t101_n_3);
  t101_g119 : ND2D0BWP7T port map(A1 => yo9, A2 => xo1, ZN => t101_n_2);
  t101_g120 : INVD0BWP7T port map(I => n_141, ZN => t101_n_1);
  t82_g136 : BUFFD4BWP7T port map(I => t82_state(1), Z => y7(12));
  t82_g141 : AN2D4BWP7T port map(A1 => t82_n_9, A2 => t82_n_10, Z => y7(13));
  t82_g185 : NR2XD0BWP7T port map(A1 => t82_n_6, A2 => reset, ZN => t82_n_8);
  t82_g186 : AOI21D0BWP7T port map(A1 => t82_n_4, A2 => t82_n_5, B => reset, ZN => t82_n_7);
  t82_g187 : AOI22D0BWP7T port map(A1 => t82_state(1), A2 => t82_n_5, B1 => t82_state(0), B2 => t82_n_3, ZN => t82_n_6);
  t82_g188 : ND3D0BWP7T port map(A1 => yo7, A2 => xo4, A3 => t82_n_2, ZN => t82_n_5);
  t82_g189 : ND2D1BWP7T port map(A1 => t82_state(0), A2 => t82_n_2, ZN => t82_n_4);
  t82_drc_bufs : INVD0BWP7T port map(I => t82_n_3, ZN => t82_n_2);
  t82_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t82_n_3);
  t82_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t82_n_7, Q => t82_state(0), QN => t82_n_10);
  t82_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t82_n_8, Q => t82_state(1), QN => t82_n_9);
  tt16_g68 : INVD4BWP7T port map(I => tt16_state, ZN => y1(12));
  tt16_state_reg : DFQD1BWP7T port map(CP => clk, D => tt16_n_3, Q => tt16_state);
  tt16_g118 : AOI211XD0BWP7T port map(A1 => y1(12), A2 => tt16_n_2, B => n_126, C => tt16_n_1, ZN => tt16_n_3);
  tt16_g119 : ND2D0BWP7T port map(A1 => xo4, A2 => yo1, ZN => tt16_n_2);
  tt16_g120 : INVD0BWP7T port map(I => lethal, ZN => tt16_n_1);
  t102_g68 : INVD4BWP7T port map(I => t102_state, ZN => y9(16));
  t102_state_reg : DFQD1BWP7T port map(CP => clk, D => t102_n_3, Q => t102_state);
  t102_g118 : AOI211XD0BWP7T port map(A1 => y9(16), A2 => t102_n_2, B => n_126, C => t102_n_1, ZN => t102_n_3);
  t102_g119 : ND2D0BWP7T port map(A1 => yo9, A2 => xo2, ZN => t102_n_2);
  t102_g120 : INVD0BWP7T port map(I => lethal, ZN => t102_n_1);
  t83_g136 : BUFFD4BWP7T port map(I => t83_state(1), Z => y7(10));
  t83_g141 : AN2D4BWP7T port map(A1 => t83_n_9, A2 => t83_n_11, Z => y7(11));
  t83_g185 : NR2XD0BWP7T port map(A1 => t83_n_6, A2 => reset, ZN => t83_n_8);
  t83_g186 : AOI21D0BWP7T port map(A1 => t83_n_4, A2 => t83_n_5, B => reset, ZN => t83_n_7);
  t83_g187 : AOI22D0BWP7T port map(A1 => t83_state(1), A2 => t83_n_5, B1 => t83_state(0), B2 => t83_n_3, ZN => t83_n_6);
  t83_g188 : ND3D0BWP7T port map(A1 => xo5, A2 => yo7, A3 => t83_n_2, ZN => t83_n_5);
  t83_g189 : ND2D1BWP7T port map(A1 => t83_state(0), A2 => t83_n_2, ZN => t83_n_4);
  t83_drc_bufs : INVD0BWP7T port map(I => t83_n_3, ZN => t83_n_2);
  t83_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t83_n_3);
  t83_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t83_n_7, Q => t83_state(0), QN => t83_n_11);
  t83_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t83_n_8, Q => t83_state(1), QN => t83_n_9);
  tt17_g68 : INVD4BWP7T port map(I => tt17_state, ZN => y1(10));
  tt17_state_reg : DFQD1BWP7T port map(CP => clk, D => tt17_n_3, Q => tt17_state);
  tt17_g118 : AOI211XD0BWP7T port map(A1 => y1(10), A2 => tt17_n_2, B => reset, C => tt17_n_1, ZN => tt17_n_3);
  tt17_g119 : ND2D0BWP7T port map(A1 => xo5, A2 => yo1, ZN => tt17_n_2);
  tt17_g120 : INVD0BWP7T port map(I => lethal, ZN => tt17_n_1);
  t103_g68 : INVD4BWP7T port map(I => t103_state, ZN => y9(14));
  t103_state_reg : DFQD1BWP7T port map(CP => clk, D => t103_n_3, Q => t103_state);
  t103_g118 : AOI211XD0BWP7T port map(A1 => y9(14), A2 => t103_n_2, B => reset, C => t103_n_1, ZN => t103_n_3);
  t103_g119 : ND2D0BWP7T port map(A1 => xo3, A2 => yo9, ZN => t103_n_2);
  t103_g120 : INVD0BWP7T port map(I => lethal, ZN => t103_n_1);
  t13_g68 : INVD4BWP7T port map(I => t13_state, ZN => y1(18));
  t13_state_reg : DFQD1BWP7T port map(CP => clk, D => t13_n_3, Q => t13_state);
  t13_g118 : AOI211XD0BWP7T port map(A1 => y1(18), A2 => t13_n_2, B => n_126, C => t13_n_1, ZN => t13_n_3);
  t13_g119 : ND2D0BWP7T port map(A1 => xo1, A2 => yo1, ZN => t13_n_2);
  t13_g120 : INVD0BWP7T port map(I => n_141, ZN => t13_n_1);
  t84_g136 : BUFFD4BWP7T port map(I => t84_state(1), Z => y7(8));
  t84_g141 : AN2D4BWP7T port map(A1 => t84_n_9, A2 => t84_n_10, Z => y7(9));
  t84_g185 : NR2XD0BWP7T port map(A1 => t84_n_6, A2 => t84_n_1, ZN => t84_n_8);
  t84_g186 : AOI21D0BWP7T port map(A1 => t84_n_4, A2 => t84_n_5, B => t84_n_1, ZN => t84_n_7);
  t84_g187 : AOI22D0BWP7T port map(A1 => t84_state(1), A2 => t84_n_5, B1 => t84_state(0), B2 => t84_n_3, ZN => t84_n_6);
  t84_g188 : ND3D0BWP7T port map(A1 => yo7, A2 => xo6, A3 => t84_n_2, ZN => t84_n_5);
  t84_g189 : ND2D1BWP7T port map(A1 => t84_state(0), A2 => t84_n_2, ZN => t84_n_4);
  t84_drc_bufs : INVD0BWP7T port map(I => t84_n_3, ZN => t84_n_2);
  t84_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t84_n_3);
  t84_drc_bufs194 : INVD0BWP7T port map(I => t84_n_0, ZN => t84_n_1);
  t84_drc_bufs196 : INVD0BWP7T port map(I => reset, ZN => t84_n_0);
  t84_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t84_n_7, Q => t84_state(0), QN => t84_n_10);
  t84_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t84_n_8, Q => t84_state(1), QN => t84_n_9);
  tt18_g68 : INVD4BWP7T port map(I => tt18_state, ZN => y1(8));
  tt18_state_reg : DFQD1BWP7T port map(CP => clk, D => tt18_n_3, Q => tt18_state);
  tt18_g118 : AOI211XD0BWP7T port map(A1 => y1(8), A2 => tt18_n_2, B => n_126, C => tt18_n_1, ZN => tt18_n_3);
  tt18_g119 : ND2D0BWP7T port map(A1 => xo6, A2 => yo1, ZN => tt18_n_2);
  tt18_g120 : INVD0BWP7T port map(I => lethal, ZN => tt18_n_1);
  t104_g136 : BUFFD4BWP7T port map(I => t104_state(1), Z => y9(12));
  t104_g141 : AN2D4BWP7T port map(A1 => t104_n_9, A2 => t104_n_11, Z => y9(13));
  t104_g185 : NR2XD0BWP7T port map(A1 => t104_n_6, A2 => n_126, ZN => t104_n_8);
  t104_g186 : AOI21D0BWP7T port map(A1 => t104_n_4, A2 => t104_n_5, B => n_126, ZN => t104_n_7);
  t104_g187 : AOI22D0BWP7T port map(A1 => t104_state(1), A2 => t104_n_5, B1 => t104_state(0), B2 => t104_n_3, ZN => t104_n_6);
  t104_g188 : ND3D0BWP7T port map(A1 => xo4, A2 => yo9, A3 => t104_n_2, ZN => t104_n_5);
  t104_g189 : ND2D1BWP7T port map(A1 => t104_state(0), A2 => t104_n_2, ZN => t104_n_4);
  t104_drc_bufs : INVD0BWP7T port map(I => t104_n_3, ZN => t104_n_2);
  t104_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t104_n_3);
  t104_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t104_n_7, Q => t104_state(0), QN => t104_n_11);
  t104_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t104_n_8, Q => t104_state(1), QN => t104_n_9);
  t14_g68 : INVD4BWP7T port map(I => t14_state, ZN => y1(16));
  t14_state_reg : DFQD1BWP7T port map(CP => clk, D => t14_n_3, Q => t14_state);
  t14_g118 : AOI211XD0BWP7T port map(A1 => y1(16), A2 => t14_n_2, B => reset, C => t14_n_1, ZN => t14_n_3);
  t14_g119 : ND2D0BWP7T port map(A1 => yo1, A2 => xo2, ZN => t14_n_2);
  t14_g120 : INVD0BWP7T port map(I => lethal, ZN => t14_n_1);
  t85_g136 : BUFFD4BWP7T port map(I => t85_state(1), Z => y7(6));
  t85_g141 : AN2D4BWP7T port map(A1 => t85_n_9, A2 => t85_n_10, Z => y7(7));
  t85_g185 : NR2XD0BWP7T port map(A1 => t85_n_6, A2 => t85_n_1, ZN => t85_n_8);
  t85_g186 : AOI21D0BWP7T port map(A1 => t85_n_4, A2 => t85_n_5, B => t85_n_1, ZN => t85_n_7);
  t85_g187 : AOI22D0BWP7T port map(A1 => t85_state(1), A2 => t85_n_5, B1 => t85_state(0), B2 => t85_n_3, ZN => t85_n_6);
  t85_g188 : ND3D0BWP7T port map(A1 => xo7, A2 => yo7, A3 => n_141, ZN => t85_n_5);
  t85_g189 : ND2D1BWP7T port map(A1 => t85_state(0), A2 => n_141, ZN => t85_n_4);
  t85_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t85_n_3);
  t85_drc_bufs194 : INVD0BWP7T port map(I => t85_n_0, ZN => t85_n_1);
  t85_drc_bufs196 : INVD0BWP7T port map(I => reset, ZN => t85_n_0);
  t85_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t85_n_7, Q => t85_state(0), QN => t85_n_10);
  t85_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t85_n_8, Q => t85_state(1), QN => t85_n_9);
  t105_g136 : BUFFD4BWP7T port map(I => t105_state(1), Z => y9(10));
  t105_g141 : AN2D4BWP7T port map(A1 => t105_n_9, A2 => t105_n_11, Z => y9(11));
  t105_g185 : NR2XD0BWP7T port map(A1 => t105_n_6, A2 => n_126, ZN => t105_n_8);
  t105_g186 : AOI21D0BWP7T port map(A1 => t105_n_4, A2 => t105_n_5, B => n_126, ZN => t105_n_7);
  t105_g187 : AOI22D0BWP7T port map(A1 => t105_state(1), A2 => t105_n_5, B1 => t105_state(0), B2 => t105_n_3, ZN => t105_n_6);
  t105_g188 : ND3D0BWP7T port map(A1 => xo5, A2 => yo9, A3 => n_141, ZN => t105_n_5);
  t105_g189 : ND2D1BWP7T port map(A1 => t105_state(0), A2 => n_141, ZN => t105_n_4);
  t105_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t105_n_3);
  t105_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t105_n_7, Q => t105_state(0), QN => t105_n_11);
  t105_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t105_n_8, Q => t105_state(1), QN => t105_n_9);
  t15_g68 : INVD4BWP7T port map(I => t15_state, ZN => y1(14));
  t15_state_reg : DFQD1BWP7T port map(CP => clk, D => t15_n_3, Q => t15_state);
  t15_g118 : AOI211XD0BWP7T port map(A1 => y1(14), A2 => t15_n_2, B => reset, C => t15_n_1, ZN => t15_n_3);
  t15_g119 : ND2D0BWP7T port map(A1 => xo3, A2 => yo1, ZN => t15_n_2);
  t15_g120 : INVD0BWP7T port map(I => lethal, ZN => t15_n_1);
  t86_g135 : BUFFD4BWP7T port map(I => t86_state(1), Z => y7(4));
  t86_g141 : AN2D4BWP7T port map(A1 => t86_n_9, A2 => t86_n_10, Z => y7(5));
  t86_g185 : NR2XD0BWP7T port map(A1 => t86_n_6, A2 => n_126, ZN => t86_n_8);
  t86_g186 : AOI21D0BWP7T port map(A1 => t86_n_4, A2 => t86_n_5, B => n_126, ZN => t86_n_7);
  t86_g187 : AOI22D0BWP7T port map(A1 => t86_state(1), A2 => t86_n_5, B1 => t86_state(0), B2 => t86_n_3, ZN => t86_n_6);
  t86_g188 : ND3D0BWP7T port map(A1 => yo7, A2 => xo8, A3 => t86_n_2, ZN => t86_n_5);
  t86_g189 : ND2D1BWP7T port map(A1 => t86_state(0), A2 => t86_n_2, ZN => t86_n_4);
  t86_drc_bufs : INVD0BWP7T port map(I => t86_n_3, ZN => t86_n_2);
  t86_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t86_n_3);
  t86_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t86_n_7, Q => t86_state(0), QN => t86_n_10);
  t86_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t86_n_8, Q => t86_state(1), QN => t86_n_9);
  t106_g136 : BUFFD4BWP7T port map(I => t106_state(1), Z => y9(8));
  t106_g141 : AN2D4BWP7T port map(A1 => t106_n_9, A2 => t106_n_10, Z => y9(9));
  t106_g185 : NR2XD0BWP7T port map(A1 => t106_n_6, A2 => t106_n_1, ZN => t106_n_8);
  t106_g186 : AOI21D0BWP7T port map(A1 => t106_n_4, A2 => t106_n_5, B => t106_n_1, ZN => t106_n_7);
  t106_g187 : AOI22D0BWP7T port map(A1 => t106_state(1), A2 => t106_n_5, B1 => t106_state(0), B2 => t106_n_3, ZN => t106_n_6);
  t106_g188 : ND3D0BWP7T port map(A1 => xo6, A2 => yo9, A3 => t106_n_2, ZN => t106_n_5);
  t106_g189 : ND2D1BWP7T port map(A1 => t106_state(0), A2 => t106_n_2, ZN => t106_n_4);
  t106_drc_bufs : INVD0BWP7T port map(I => t106_n_3, ZN => t106_n_2);
  t106_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t106_n_3);
  t106_drc_bufs194 : INVD0BWP7T port map(I => t106_n_0, ZN => t106_n_1);
  t106_drc_bufs196 : INVD0BWP7T port map(I => reset, ZN => t106_n_0);
  t106_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t106_n_7, Q => t106_state(0), QN => t106_n_10);
  t106_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t106_n_8, Q => t106_state(1), QN => t106_n_9);
  t87_g68 : INVD4BWP7T port map(I => t87_state, ZN => y7(2));
  t87_state_reg : DFQD1BWP7T port map(CP => clk, D => t87_n_3, Q => t87_state);
  t87_g118 : AOI211XD0BWP7T port map(A1 => y7(2), A2 => t87_n_2, B => reset, C => t87_n_1, ZN => t87_n_3);
  t87_g119 : ND2D0BWP7T port map(A1 => yo7, A2 => xo9, ZN => t87_n_2);
  t87_g120 : INVD0BWP7T port map(I => lethal, ZN => t87_n_1);
  t107_g68 : INVD4BWP7T port map(I => t107_state, ZN => y9(6));
  t107_state_reg : DFQD1BWP7T port map(CP => clk, D => t107_n_3, Q => t107_state);
  t107_g118 : AOI211XD0BWP7T port map(A1 => y9(6), A2 => t107_n_2, B => reset, C => t107_n_1, ZN => t107_n_3);
  t107_g119 : ND2D0BWP7T port map(A1 => xo7, A2 => yo9, ZN => t107_n_2);
  t107_g120 : INVD0BWP7T port map(I => lethal, ZN => t107_n_1);
  t108_g68 : INVD4BWP7T port map(I => t108_state, ZN => y9(4));
  t108_state_reg : DFQD1BWP7T port map(CP => clk, D => t108_n_3, Q => t108_state);
  t108_g118 : AOI211XD0BWP7T port map(A1 => y9(4), A2 => t108_n_2, B => reset, C => t108_n_1, ZN => t108_n_3);
  t108_g119 : ND2D0BWP7T port map(A1 => yo9, A2 => xo8, ZN => t108_n_2);
  t108_g120 : INVD0BWP7T port map(I => lethal, ZN => t108_n_1);
  t90_g68 : INVD4BWP7T port map(I => t90_state, ZN => y8(18));
  t90_state_reg : DFQD1BWP7T port map(CP => clk, D => t90_n_3, Q => t90_state);
  t90_g118 : AOI211XD0BWP7T port map(A1 => y8(18), A2 => t90_n_2, B => reset, C => t90_n_1, ZN => t90_n_3);
  t90_g119 : ND2D0BWP7T port map(A1 => yo8, A2 => xo1, ZN => t90_n_2);
  t90_g120 : INVD0BWP7T port map(I => lethal, ZN => t90_n_1);
  t109_g68 : INVD4BWP7T port map(I => t109_state, ZN => y9(2));
  t109_state_reg : DFQD1BWP7T port map(CP => clk, D => t109_n_3, Q => t109_state);
  t109_g118 : AOI211XD0BWP7T port map(A1 => y9(2), A2 => t109_n_2, B => n_126, C => t109_n_1, ZN => t109_n_3);
  t109_g119 : ND2D0BWP7T port map(A1 => yo9, A2 => xo9, ZN => t109_n_2);
  t109_g120 : INVD0BWP7T port map(I => n_141, ZN => t109_n_1);
  t20_g68 : INVD4BWP7T port map(I => t20_state, ZN => y1(4));
  t20_state_reg : DFQD1BWP7T port map(CP => clk, D => t20_n_3, Q => t20_state);
  t20_g118 : AOI211XD0BWP7T port map(A1 => y1(4), A2 => t20_n_2, B => n_126, C => t20_n_1, ZN => t20_n_3);
  t20_g119 : ND2D0BWP7T port map(A1 => xo8, A2 => yo1, ZN => t20_n_2);
  t20_g120 : INVD0BWP7T port map(I => lethal, ZN => t20_n_1);
  t19_g68 : INVD4BWP7T port map(I => t19_state, ZN => y1(6));
  t19_state_reg : DFQD1BWP7T port map(CP => clk, D => t19_n_3, Q => t19_state);
  t19_g118 : AOI211XD0BWP7T port map(A1 => y1(6), A2 => t19_n_2, B => reset, C => t19_n_1, ZN => t19_n_3);
  t19_g119 : ND2D0BWP7T port map(A1 => xo7, A2 => yo1, ZN => t19_n_2);
  t19_g120 : INVD0BWP7T port map(I => lethal, ZN => t19_n_1);
  xyconv_g492 : INR2XD0BWP7T port map(A1 => lethalx(1), B1 => xyconv_n_16, ZN => xo7);
  xyconv_g493 : NR2XD0BWP7T port map(A1 => xyconv_n_16, A2 => lethalx(1), ZN => xo5);
  xyconv_g494 : INR2XD0BWP7T port map(A1 => lethalx(1), B1 => xyconv_n_10, ZN => xo6);
  xyconv_g495 : NR2XD0BWP7T port map(A1 => xyconv_n_11, A2 => lethaly(1), ZN => yo4);
  xyconv_g496 : NR2XD0BWP7T port map(A1 => xyconv_n_10, A2 => lethalx(1), ZN => xo4);
  xyconv_g497 : NR2XD0BWP7T port map(A1 => xyconv_n_12, A2 => lethaly(1), ZN => yo5);
  xyconv_g498 : INR2XD0BWP7T port map(A1 => lethaly(1), B1 => xyconv_n_11, ZN => yo6);
  xyconv_g499 : NR2XD0BWP7T port map(A1 => xyconv_n_15, A2 => lethalx(0), ZN => xo8);
  xyconv_g500 : NR3D0BWP7T port map(A1 => xyconv_n_3, A2 => lethaly(2), A3 => xyconv_n_1, ZN => yo3);
  xyconv_g501 : NR2XD0BWP7T port map(A1 => xyconv_n_14, A2 => lethaly(0), ZN => yo8);
  xyconv_g502 : INR2XD0BWP7T port map(A1 => lethaly(0), B1 => xyconv_n_14, ZN => yo9);
  xyconv_g503 : INR2XD0BWP7T port map(A1 => lethalx(0), B1 => xyconv_n_15, ZN => xo9);
  xyconv_g504 : INR2XD0BWP7T port map(A1 => lethaly(1), B1 => xyconv_n_12, ZN => yo7);
  xyconv_g505 : NR3D0BWP7T port map(A1 => xyconv_n_6, A2 => lethalx(2), A3 => xyconv_n_2, ZN => xo2);
  xyconv_g506 : NR3D0BWP7T port map(A1 => xyconv_n_4, A2 => lethalx(2), A3 => xyconv_n_2, ZN => xo3);
  xyconv_g507 : NR3D0BWP7T port map(A1 => xyconv_n_8, A2 => lethaly(2), A3 => xyconv_n_1, ZN => yo2);
  xyconv_g508 : INR2XD0BWP7T port map(A1 => xyconv_n_5, B1 => xyconv_n_4, ZN => xo1);
  xyconv_g509 : IND2D1BWP7T port map(A1 => xyconv_n_4, B1 => lethalx(2), ZN => xyconv_n_16);
  xyconv_g510 : ND2D1BWP7T port map(A1 => xyconv_n_5, A2 => lethalx(3), ZN => xyconv_n_15);
  xyconv_g511 : ND2D1BWP7T port map(A1 => xyconv_n_7, A2 => lethaly(3), ZN => xyconv_n_14);
  xyconv_g512 : INR2XD0BWP7T port map(A1 => xyconv_n_7, B1 => xyconv_n_3, ZN => yo1);
  xyconv_g513 : IND2D1BWP7T port map(A1 => xyconv_n_3, B1 => lethaly(2), ZN => xyconv_n_12);
  xyconv_g514 : IND2D1BWP7T port map(A1 => xyconv_n_8, B1 => lethaly(2), ZN => xyconv_n_11);
  xyconv_g515 : IND2D1BWP7T port map(A1 => xyconv_n_6, B1 => lethalx(2), ZN => xyconv_n_10);
  xyconv_g516 : OR2D1BWP7T port map(A1 => lethaly(3), A2 => lethaly(0), Z => xyconv_n_8);
  xyconv_g517 : NR2XD0BWP7T port map(A1 => lethaly(1), A2 => lethaly(2), ZN => xyconv_n_7);
  xyconv_g518 : OR2D1BWP7T port map(A1 => lethalx(3), A2 => lethalx(0), Z => xyconv_n_6);
  xyconv_g519 : NR2XD0BWP7T port map(A1 => lethalx(1), A2 => lethalx(2), ZN => xyconv_n_5);
  xyconv_g520 : IND2D1BWP7T port map(A1 => lethalx(3), B1 => lethalx(0), ZN => xyconv_n_4);
  xyconv_g521 : IND2D1BWP7T port map(A1 => lethaly(3), B1 => lethaly(0), ZN => xyconv_n_3);
  xyconv_g522 : INVD1BWP7T port map(I => lethalx(1), ZN => xyconv_n_2);
  xyconv_g523 : INVD1BWP7T port map(I => lethaly(1), ZN => xyconv_n_1);
  t92_g135 : BUFFD4BWP7T port map(I => t92_state(1), Z => y8(14));
  t92_g141 : AN2D4BWP7T port map(A1 => t92_n_9, A2 => t92_n_11, Z => y8(15));
  t92_g185 : NR2XD0BWP7T port map(A1 => t92_n_6, A2 => n_126, ZN => t92_n_8);
  t92_g186 : AOI21D0BWP7T port map(A1 => t92_n_4, A2 => t92_n_5, B => n_126, ZN => t92_n_7);
  t92_g187 : AOI22D0BWP7T port map(A1 => t92_state(1), A2 => t92_n_5, B1 => t92_state(0), B2 => t92_n_3, ZN => t92_n_6);
  t92_g188 : ND3D0BWP7T port map(A1 => xo3, A2 => yo8, A3 => n_141, ZN => t92_n_5);
  t92_g189 : ND2D1BWP7T port map(A1 => t92_state(0), A2 => n_141, ZN => t92_n_4);
  t92_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t92_n_3);
  t92_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t92_n_7, Q => t92_state(0), QN => t92_n_11);
  t92_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t92_n_8, Q => t92_state(1), QN => t92_n_9);
  t21_g68 : INVD4BWP7T port map(I => t21_state, ZN => y1(2));
  t21_state_reg : DFQD1BWP7T port map(CP => clk, D => t21_n_3, Q => t21_state);
  t21_g118 : AOI211XD0BWP7T port map(A1 => y1(2), A2 => t21_n_2, B => n_126, C => t21_n_1, ZN => t21_n_3);
  t21_g119 : ND2D0BWP7T port map(A1 => xo9, A2 => yo1, ZN => t21_n_2);
  t21_g120 : INVD0BWP7T port map(I => n_141, ZN => t21_n_1);
  t94_g136 : BUFFD4BWP7T port map(I => t94_state(1), Z => y8(10));
  t94_g141 : AN2D4BWP7T port map(A1 => t94_n_9, A2 => t94_n_10, Z => y8(11));
  t94_g185 : NR2XD0BWP7T port map(A1 => t94_n_6, A2 => reset, ZN => t94_n_8);
  t94_g186 : AOI21D0BWP7T port map(A1 => t94_n_4, A2 => t94_n_5, B => reset, ZN => t94_n_7);
  t94_g187 : AOI22D0BWP7T port map(A1 => t94_state(1), A2 => t94_n_5, B1 => t94_state(0), B2 => t94_n_3, ZN => t94_n_6);
  t94_g188 : ND3D0BWP7T port map(A1 => xo5, A2 => yo8, A3 => t94_n_2, ZN => t94_n_5);
  t94_g189 : ND2D1BWP7T port map(A1 => t94_state(0), A2 => t94_n_2, ZN => t94_n_4);
  t94_drc_bufs : INVD0BWP7T port map(I => t94_n_3, ZN => t94_n_2);
  t94_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t94_n_3);
  t94_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t94_n_7, Q => t94_state(0), QN => t94_n_10);
  t94_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t94_n_8, Q => t94_state(1), QN => t94_n_9);
  t24_g68 : INVD4BWP7T port map(I => t24_state, ZN => y2(18));
  t24_state_reg : DFQD1BWP7T port map(CP => clk, D => t24_n_3, Q => t24_state);
  t24_g118 : AOI211XD0BWP7T port map(A1 => y2(18), A2 => t24_n_2, B => n_126, C => t24_n_1, ZN => t24_n_3);
  t24_g119 : ND2D0BWP7T port map(A1 => xo1, A2 => yo2, ZN => t24_n_2);
  t24_g120 : INVD0BWP7T port map(I => lethal, ZN => t24_n_1);
  t96_g136 : BUFFD4BWP7T port map(I => t96_state(1), Z => y8(6));
  t96_g141 : AN2D4BWP7T port map(A1 => t96_n_9, A2 => t96_n_11, Z => y8(7));
  t96_g185 : NR2XD0BWP7T port map(A1 => t96_n_6, A2 => reset, ZN => t96_n_8);
  t96_g186 : AOI21D0BWP7T port map(A1 => t96_n_4, A2 => t96_n_5, B => reset, ZN => t96_n_7);
  t96_g187 : AOI22D0BWP7T port map(A1 => t96_state(1), A2 => t96_n_5, B1 => t96_state(0), B2 => t96_n_3, ZN => t96_n_6);
  t96_g188 : ND3D0BWP7T port map(A1 => xo7, A2 => yo8, A3 => t96_n_2, ZN => t96_n_5);
  t96_g189 : ND2D1BWP7T port map(A1 => t96_state(0), A2 => t96_n_2, ZN => t96_n_4);
  t96_drc_bufs : INVD0BWP7T port map(I => t96_n_3, ZN => t96_n_2);
  t96_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t96_n_3);
  t96_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t96_n_7, Q => t96_state(0), QN => t96_n_11);
  t96_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t96_n_8, Q => t96_state(1), QN => t96_n_9);
  t26_g136 : BUFFD4BWP7T port map(I => t26_state(1), Z => y2(14));
  t26_g141 : AN2D4BWP7T port map(A1 => t26_n_9, A2 => t26_n_10, Z => y2(15));
  t26_g185 : NR2XD0BWP7T port map(A1 => t26_n_6, A2 => reset, ZN => t26_n_8);
  t26_g186 : AOI21D0BWP7T port map(A1 => t26_n_4, A2 => t26_n_5, B => reset, ZN => t26_n_7);
  t26_g187 : AOI22D0BWP7T port map(A1 => t26_state(1), A2 => t26_n_5, B1 => t26_state(0), B2 => t26_n_3, ZN => t26_n_6);
  t26_g188 : ND3D0BWP7T port map(A1 => xo3, A2 => yo2, A3 => t26_n_2, ZN => t26_n_5);
  t26_g189 : ND2D1BWP7T port map(A1 => t26_state(0), A2 => t26_n_2, ZN => t26_n_4);
  t26_drc_bufs : INVD0BWP7T port map(I => t26_n_3, ZN => t26_n_2);
  t26_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t26_n_3);
  t26_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t26_n_7, Q => t26_state(0), QN => t26_n_10);
  t26_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t26_n_8, Q => t26_state(1), QN => t26_n_9);
  t98_g68 : INVD4BWP7T port map(I => t98_state, ZN => y8(2));
  t98_state_reg : DFQD1BWP7T port map(CP => clk, D => t98_n_3, Q => t98_state);
  t98_g118 : AOI211XD0BWP7T port map(A1 => y8(2), A2 => t98_n_2, B => reset, C => t98_n_1, ZN => t98_n_3);
  t98_g119 : ND2D0BWP7T port map(A1 => xo9, A2 => yo8, ZN => t98_n_2);
  t98_g120 : INVD0BWP7T port map(I => lethal, ZN => t98_n_1);
  t28_g136 : BUFFD4BWP7T port map(I => t28_state(1), Z => y2(10));
  t28_g141 : AN2D4BWP7T port map(A1 => t28_n_9, A2 => t28_n_10, Z => y2(11));
  t28_g185 : NR2XD0BWP7T port map(A1 => t28_n_6, A2 => n_126, ZN => t28_n_8);
  t28_g186 : AOI21D0BWP7T port map(A1 => t28_n_4, A2 => t28_n_5, B => n_126, ZN => t28_n_7);
  t28_g187 : AOI22D0BWP7T port map(A1 => t28_state(1), A2 => t28_n_5, B1 => t28_state(0), B2 => t28_n_3, ZN => t28_n_6);
  t28_g188 : ND3D0BWP7T port map(A1 => xo5, A2 => yo2, A3 => t28_n_2, ZN => t28_n_5);
  t28_g189 : ND2D1BWP7T port map(A1 => t28_state(0), A2 => t28_n_2, ZN => t28_n_4);
  t28_drc_bufs : INVD0BWP7T port map(I => t28_n_3, ZN => t28_n_2);
  t28_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t28_n_3);
  t28_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t28_n_7, Q => t28_state(0), QN => t28_n_10);
  t28_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t28_n_8, Q => t28_state(1), QN => t28_n_9);
  t30_g136 : BUFFD4BWP7T port map(I => t30_state(1), Z => y2(6));
  t30_g141 : AN2D4BWP7T port map(A1 => t30_n_9, A2 => t30_n_10, Z => y2(7));
  t30_g185 : NR2XD0BWP7T port map(A1 => t30_n_6, A2 => n_126, ZN => t30_n_8);
  t30_g186 : AOI21D0BWP7T port map(A1 => t30_n_4, A2 => t30_n_5, B => n_126, ZN => t30_n_7);
  t30_g187 : AOI22D0BWP7T port map(A1 => t30_state(1), A2 => t30_n_5, B1 => t30_state(0), B2 => t30_n_3, ZN => t30_n_6);
  t30_g188 : ND3D0BWP7T port map(A1 => xo7, A2 => yo2, A3 => n_141, ZN => t30_n_5);
  t30_g189 : ND2D1BWP7T port map(A1 => t30_state(0), A2 => n_141, ZN => t30_n_4);
  t30_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t30_n_3);
  t30_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t30_n_7, Q => t30_state(0), QN => t30_n_10);
  t30_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t30_n_8, Q => t30_state(1), QN => t30_n_9);
  t32_g68 : INVD4BWP7T port map(I => t32_state, ZN => y2(2));
  t32_state_reg : DFQD1BWP7T port map(CP => clk, D => t32_n_3, Q => t32_state);
  t32_g118 : AOI211XD0BWP7T port map(A1 => y2(2), A2 => t32_n_2, B => n_126, C => t32_n_1, ZN => t32_n_3);
  t32_g119 : ND2D0BWP7T port map(A1 => xo9, A2 => yo2, ZN => t32_n_2);
  t32_g120 : INVD0BWP7T port map(I => lethal, ZN => t32_n_1);
  t35_g68 : INVD4BWP7T port map(I => t35_state, ZN => y3(18));
  t35_state_reg : DFQD1BWP7T port map(CP => clk, D => t35_n_3, Q => t35_state);
  t35_g118 : AOI211XD0BWP7T port map(A1 => y3(18), A2 => t35_n_2, B => reset, C => t35_n_1, ZN => t35_n_3);
  t35_g119 : ND2D0BWP7T port map(A1 => yo3, A2 => xo1, ZN => t35_n_2);
  t35_g120 : INVD0BWP7T port map(I => lethal, ZN => t35_n_1);
  t36_g136 : BUFFD4BWP7T port map(I => t36_state(1), Z => y3(16));
  t36_g141 : AN2D4BWP7T port map(A1 => t36_n_9, A2 => t36_n_10, Z => y3(17));
  t36_g185 : NR2XD0BWP7T port map(A1 => t36_n_6, A2 => n_126, ZN => t36_n_8);
  t36_g186 : AOI21D0BWP7T port map(A1 => t36_n_4, A2 => t36_n_5, B => n_126, ZN => t36_n_7);
  t36_g187 : AOI22D0BWP7T port map(A1 => t36_state(1), A2 => t36_n_5, B1 => t36_state(0), B2 => t36_n_3, ZN => t36_n_6);
  t36_g188 : ND3D0BWP7T port map(A1 => yo3, A2 => xo2, A3 => t36_n_2, ZN => t36_n_5);
  t36_g189 : ND2D1BWP7T port map(A1 => t36_state(0), A2 => t36_n_2, ZN => t36_n_4);
  t36_drc_bufs : INVD0BWP7T port map(I => t36_n_3, ZN => t36_n_2);
  t36_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t36_n_3);
  t36_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t36_n_7, Q => t36_state(0), QN => t36_n_10);
  t36_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t36_n_8, Q => t36_state(1), QN => t36_n_9);
  t37_g136 : BUFFD4BWP7T port map(I => t37_state(1), Z => y3(14));
  t37_g141 : AN2D4BWP7T port map(A1 => t37_n_9, A2 => t37_n_10, Z => y3(15));
  t37_g185 : NR2XD0BWP7T port map(A1 => t37_n_6, A2 => n_126, ZN => t37_n_8);
  t37_g186 : AOI21D0BWP7T port map(A1 => t37_n_4, A2 => t37_n_5, B => n_126, ZN => t37_n_7);
  t37_g187 : AOI22D0BWP7T port map(A1 => t37_state(1), A2 => t37_n_5, B1 => t37_state(0), B2 => t37_n_3, ZN => t37_n_6);
  t37_g188 : ND3D0BWP7T port map(A1 => xo3, A2 => yo3, A3 => n_141, ZN => t37_n_5);
  t37_g189 : ND2D1BWP7T port map(A1 => t37_state(0), A2 => n_141, ZN => t37_n_4);
  t37_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t37_n_3);
  t37_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t37_n_7, Q => t37_state(0), QN => t37_n_10);
  t37_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t37_n_8, Q => t37_state(1), QN => t37_n_9);
  t38_g135 : BUFFD4BWP7T port map(I => t38_state(1), Z => y3(12));
  t38_g141 : AN2D4BWP7T port map(A1 => t38_n_9, A2 => t38_n_10, Z => y3(13));
  t38_g185 : NR2XD0BWP7T port map(A1 => t38_n_6, A2 => reset, ZN => t38_n_8);
  t38_g186 : AOI21D0BWP7T port map(A1 => t38_n_4, A2 => t38_n_5, B => reset, ZN => t38_n_7);
  t38_g187 : AOI22D0BWP7T port map(A1 => t38_state(1), A2 => t38_n_5, B1 => t38_state(0), B2 => t38_n_3, ZN => t38_n_6);
  t38_g188 : ND3D0BWP7T port map(A1 => yo3, A2 => xo4, A3 => t38_n_2, ZN => t38_n_5);
  t38_g189 : ND2D1BWP7T port map(A1 => t38_state(0), A2 => t38_n_2, ZN => t38_n_4);
  t38_drc_bufs : INVD0BWP7T port map(I => t38_n_3, ZN => t38_n_2);
  t38_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t38_n_3);
  t38_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t38_n_7, Q => t38_state(0), QN => t38_n_10);
  t38_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t38_n_8, Q => t38_state(1), QN => t38_n_9);
  t39_g135 : BUFFD4BWP7T port map(I => t39_state(1), Z => y3(10));
  t39_g141 : AN2D4BWP7T port map(A1 => t39_n_9, A2 => t39_n_10, Z => y3(11));
  t39_g185 : NR2XD0BWP7T port map(A1 => t39_n_6, A2 => t39_n_1, ZN => t39_n_8);
  t39_g186 : AOI21D0BWP7T port map(A1 => t39_n_4, A2 => t39_n_5, B => t39_n_1, ZN => t39_n_7);
  t39_g187 : AOI22D0BWP7T port map(A1 => t39_state(1), A2 => t39_n_5, B1 => t39_state(0), B2 => t39_n_3, ZN => t39_n_6);
  t39_g188 : ND3D0BWP7T port map(A1 => xo5, A2 => yo3, A3 => t39_n_2, ZN => t39_n_5);
  t39_g189 : ND2D1BWP7T port map(A1 => t39_state(0), A2 => t39_n_2, ZN => t39_n_4);
  t39_drc_bufs : INVD0BWP7T port map(I => t39_n_3, ZN => t39_n_2);
  t39_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t39_n_3);
  t39_drc_bufs194 : INVD0BWP7T port map(I => t39_n_0, ZN => t39_n_1);
  t39_drc_bufs196 : INVD0BWP7T port map(I => reset, ZN => t39_n_0);
  t39_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t39_n_7, Q => t39_state(0), QN => t39_n_10);
  t39_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t39_n_8, Q => t39_state(1), QN => t39_n_9);
  t40_g136 : BUFFD4BWP7T port map(I => t40_state(1), Z => y3(8));
  t40_g141 : AN2D4BWP7T port map(A1 => t40_n_9, A2 => t40_n_10, Z => y3(9));
  t40_g185 : NR2XD0BWP7T port map(A1 => t40_n_6, A2 => n_126, ZN => t40_n_8);
  t40_g186 : AOI21D0BWP7T port map(A1 => t40_n_4, A2 => t40_n_5, B => n_126, ZN => t40_n_7);
  t40_g187 : AOI22D0BWP7T port map(A1 => t40_state(1), A2 => t40_n_5, B1 => t40_state(0), B2 => t40_n_3, ZN => t40_n_6);
  t40_g188 : ND3D0BWP7T port map(A1 => yo3, A2 => xo6, A3 => t40_n_2, ZN => t40_n_5);
  t40_g189 : ND2D1BWP7T port map(A1 => t40_state(0), A2 => t40_n_2, ZN => t40_n_4);
  t40_drc_bufs : INVD0BWP7T port map(I => t40_n_3, ZN => t40_n_2);
  t40_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t40_n_3);
  t40_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t40_n_7, Q => t40_state(0), QN => t40_n_10);
  t40_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t40_n_8, Q => t40_state(1), QN => t40_n_9);
  t41_g136 : BUFFD4BWP7T port map(I => t41_state(1), Z => y3(6));
  t41_g141 : AN2D4BWP7T port map(A1 => t41_n_9, A2 => t41_n_10, Z => y3(7));
  t41_g185 : NR2XD0BWP7T port map(A1 => t41_n_6, A2 => n_126, ZN => t41_n_8);
  t41_g186 : AOI21D0BWP7T port map(A1 => t41_n_4, A2 => t41_n_5, B => n_126, ZN => t41_n_7);
  t41_g187 : AOI22D0BWP7T port map(A1 => t41_state(1), A2 => t41_n_5, B1 => t41_state(0), B2 => t41_n_3, ZN => t41_n_6);
  t41_g188 : ND3D0BWP7T port map(A1 => xo7, A2 => yo3, A3 => n_141, ZN => t41_n_5);
  t41_g189 : ND2D1BWP7T port map(A1 => t41_state(0), A2 => n_141, ZN => t41_n_4);
  t41_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t41_n_3);
  t41_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t41_n_7, Q => t41_state(0), QN => t41_n_10);
  t41_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t41_n_8, Q => t41_state(1), QN => t41_n_9);
  t42_g135 : BUFFD4BWP7T port map(I => t42_state(1), Z => y3(4));
  t42_g141 : AN2D4BWP7T port map(A1 => t42_n_9, A2 => t42_n_10, Z => y3(5));
  t42_g185 : NR2XD0BWP7T port map(A1 => t42_n_6, A2 => t42_n_1, ZN => t42_n_8);
  t42_g186 : AOI21D0BWP7T port map(A1 => t42_n_4, A2 => t42_n_5, B => t42_n_1, ZN => t42_n_7);
  t42_g187 : AOI22D0BWP7T port map(A1 => t42_state(1), A2 => t42_n_5, B1 => t42_state(0), B2 => t42_n_3, ZN => t42_n_6);
  t42_g188 : ND3D0BWP7T port map(A1 => yo3, A2 => xo8, A3 => t42_n_2, ZN => t42_n_5);
  t42_g189 : ND2D1BWP7T port map(A1 => t42_state(0), A2 => t42_n_2, ZN => t42_n_4);
  t42_drc_bufs : INVD0BWP7T port map(I => t42_n_3, ZN => t42_n_2);
  t42_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t42_n_3);
  t42_drc_bufs194 : INVD0BWP7T port map(I => t42_n_0, ZN => t42_n_1);
  t42_drc_bufs196 : INVD0BWP7T port map(I => reset, ZN => t42_n_0);
  t42_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t42_n_7, Q => t42_state(0), QN => t42_n_10);
  t42_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t42_n_8, Q => t42_state(1), QN => t42_n_9);
  t43_g68 : INVD4BWP7T port map(I => t43_state, ZN => y3(2));
  t43_state_reg : DFQD1BWP7T port map(CP => clk, D => t43_n_3, Q => t43_state);
  t43_g118 : AOI211XD0BWP7T port map(A1 => y3(2), A2 => t43_n_2, B => reset, C => t43_n_1, ZN => t43_n_3);
  t43_g119 : ND2D0BWP7T port map(A1 => yo3, A2 => xo9, ZN => t43_n_2);
  t43_g120 : INVD0BWP7T port map(I => lethal, ZN => t43_n_1);
  t46_g135 : BUFFD4BWP7T port map(I => t46_state(1), Z => y4(18));
  t46_g141 : AN2D4BWP7T port map(A1 => t46_n_9, A2 => t46_n_11, Z => y4(19));
  t46_g185 : NR2XD0BWP7T port map(A1 => t46_n_6, A2 => n_126, ZN => t46_n_8);
  t46_g186 : AOI21D0BWP7T port map(A1 => t46_n_4, A2 => t46_n_5, B => n_126, ZN => t46_n_7);
  t46_g187 : AOI22D0BWP7T port map(A1 => t46_state(1), A2 => t46_n_5, B1 => t46_state(0), B2 => t46_n_3, ZN => t46_n_6);
  t46_g188 : ND3D0BWP7T port map(A1 => yo4, A2 => xo1, A3 => t46_n_2, ZN => t46_n_5);
  t46_g189 : ND2D1BWP7T port map(A1 => t46_state(0), A2 => t46_n_2, ZN => t46_n_4);
  t46_drc_bufs : INVD0BWP7T port map(I => t46_n_3, ZN => t46_n_2);
  t46_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t46_n_3);
  t46_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t46_n_7, Q => t46_state(0), QN => t46_n_11);
  t46_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t46_n_8, Q => t46_state(1), QN => t46_n_9);
  t48_g136 : BUFFD4BWP7T port map(I => t48_state(1), Z => y4(14));
  t48_g141 : AN2D4BWP7T port map(A1 => t48_n_9, A2 => t48_n_10, Z => y4(15));
  t48_g185 : NR2XD0BWP7T port map(A1 => t48_n_6, A2 => n_126, ZN => t48_n_8);
  t48_g186 : AOI21D0BWP7T port map(A1 => t48_n_4, A2 => t48_n_5, B => n_126, ZN => t48_n_7);
  t48_g187 : AOI22D0BWP7T port map(A1 => t48_state(1), A2 => t48_n_5, B1 => t48_state(0), B2 => t48_n_3, ZN => t48_n_6);
  t48_g188 : ND3D0BWP7T port map(A1 => xo3, A2 => yo4, A3 => n_141, ZN => t48_n_5);
  t48_g189 : ND2D1BWP7T port map(A1 => t48_state(0), A2 => n_141, ZN => t48_n_4);
  t48_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t48_n_3);
  t48_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t48_n_7, Q => t48_state(0), QN => t48_n_10);
  t48_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t48_n_8, Q => t48_state(1), QN => t48_n_9);
  t50_g68 : INVD4BWP7T port map(I => t50_state, ZN => y4(10));
  t50_state_reg : DFQD1BWP7T port map(CP => clk, D => t50_n_3, Q => t50_state);
  t50_g118 : AOI211XD0BWP7T port map(A1 => y4(10), A2 => t50_n_2, B => n_126, C => t50_n_1, ZN => t50_n_3);
  t50_g119 : ND2D0BWP7T port map(A1 => xo5, A2 => yo4, ZN => t50_n_2);
  t50_g120 : INVD0BWP7T port map(I => lethal, ZN => t50_n_1);
  t52_g136 : BUFFD4BWP7T port map(I => t52_state(1), Z => y4(6));
  t52_g141 : AN2D4BWP7T port map(A1 => t52_n_9, A2 => t52_n_11, Z => y4(7));
  t52_g185 : NR2XD0BWP7T port map(A1 => t52_n_6, A2 => t52_n_1, ZN => t52_n_8);
  t52_g186 : AOI21D0BWP7T port map(A1 => t52_n_4, A2 => t52_n_5, B => t52_n_1, ZN => t52_n_7);
  t52_g187 : AOI22D0BWP7T port map(A1 => t52_state(1), A2 => t52_n_5, B1 => t52_state(0), B2 => t52_n_3, ZN => t52_n_6);
  t52_g188 : ND3D0BWP7T port map(A1 => xo7, A2 => yo4, A3 => t52_n_2, ZN => t52_n_5);
  t52_g189 : ND2D1BWP7T port map(A1 => t52_state(0), A2 => t52_n_2, ZN => t52_n_4);
  t52_drc_bufs : INVD0BWP7T port map(I => t52_n_3, ZN => t52_n_2);
  t52_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t52_n_3);
  t52_drc_bufs194 : INVD0BWP7T port map(I => t52_n_0, ZN => t52_n_1);
  t52_drc_bufs196 : INVD0BWP7T port map(I => reset, ZN => t52_n_0);
  t52_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t52_n_7, Q => t52_state(0), QN => t52_n_11);
  t52_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t52_n_8, Q => t52_state(1), QN => t52_n_9);
  t54_g135 : BUFFD4BWP7T port map(I => t54_state(1), Z => y4(2));
  t54_g141 : AN2D4BWP7T port map(A1 => t54_n_9, A2 => t54_n_11, Z => y4(3));
  t54_g185 : NR2XD0BWP7T port map(A1 => t54_n_6, A2 => n_126, ZN => t54_n_8);
  t54_g186 : AOI21D0BWP7T port map(A1 => t54_n_4, A2 => t54_n_5, B => n_126, ZN => t54_n_7);
  t54_g187 : AOI22D0BWP7T port map(A1 => t54_state(1), A2 => t54_n_5, B1 => t54_state(0), B2 => t54_n_3, ZN => t54_n_6);
  t54_g188 : ND3D0BWP7T port map(A1 => yo4, A2 => xo9, A3 => t54_n_2, ZN => t54_n_5);
  t54_g189 : ND2D1BWP7T port map(A1 => t54_state(0), A2 => t54_n_2, ZN => t54_n_4);
  t54_drc_bufs : INVD0BWP7T port map(I => t54_n_3, ZN => t54_n_2);
  t54_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t54_n_3);
  t54_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t54_n_7, Q => t54_state(0), QN => t54_n_11);
  t54_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t54_n_8, Q => t54_state(1), QN => t54_n_9);
  t57_g136 : BUFFD4BWP7T port map(I => t57_state(1), Z => y5(18));
  t57_g141 : AN2D4BWP7T port map(A1 => t57_n_9, A2 => t57_n_11, Z => y5(19));
  t57_g185 : NR2XD0BWP7T port map(A1 => t57_n_6, A2 => n_126, ZN => t57_n_8);
  t57_g186 : AOI21D0BWP7T port map(A1 => t57_n_4, A2 => t57_n_5, B => n_126, ZN => t57_n_7);
  t57_g187 : AOI22D0BWP7T port map(A1 => t57_state(1), A2 => t57_n_5, B1 => t57_state(0), B2 => t57_n_3, ZN => t57_n_6);
  t57_g188 : ND3D0BWP7T port map(A1 => yo5, A2 => xo1, A3 => n_141, ZN => t57_n_5);
  t57_g189 : ND2D1BWP7T port map(A1 => t57_state(0), A2 => n_141, ZN => t57_n_4);
  t57_drc_bufs192 : INVD0BWP7T port map(I => n_141, ZN => t57_n_3);
  t57_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t57_n_7, Q => t57_state(0), QN => t57_n_11);
  t57_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t57_n_8, Q => t57_state(1), QN => t57_n_9);
  t58_g136 : BUFFD4BWP7T port map(I => t58_state(1), Z => y5(16));
  t58_g141 : AN2D4BWP7T port map(A1 => t58_n_9, A2 => t58_n_10, Z => y5(17));
  t58_g185 : NR2XD0BWP7T port map(A1 => t58_n_6, A2 => t58_n_1, ZN => t58_n_8);
  t58_g186 : AOI21D0BWP7T port map(A1 => t58_n_4, A2 => t58_n_5, B => t58_n_1, ZN => t58_n_7);
  t58_g187 : AOI22D0BWP7T port map(A1 => t58_state(1), A2 => t58_n_5, B1 => t58_state(0), B2 => t58_n_3, ZN => t58_n_6);
  t58_g188 : ND3D0BWP7T port map(A1 => yo5, A2 => xo2, A3 => t58_n_2, ZN => t58_n_5);
  t58_g189 : ND2D1BWP7T port map(A1 => t58_state(0), A2 => t58_n_2, ZN => t58_n_4);
  t58_drc_bufs : INVD0BWP7T port map(I => t58_n_3, ZN => t58_n_2);
  t58_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t58_n_3);
  t58_drc_bufs194 : INVD0BWP7T port map(I => t58_n_0, ZN => t58_n_1);
  t58_drc_bufs196 : INVD0BWP7T port map(I => reset, ZN => t58_n_0);
  t58_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t58_n_7, Q => t58_state(0), QN => t58_n_10);
  t58_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t58_n_8, Q => t58_state(1), QN => t58_n_9);
  t59_g136 : BUFFD4BWP7T port map(I => t59_state(1), Z => y5(14));
  t59_g141 : AN2D4BWP7T port map(A1 => t59_n_9, A2 => t59_n_11, Z => y5(15));
  t59_g185 : NR2XD0BWP7T port map(A1 => t59_n_6, A2 => reset, ZN => t59_n_8);
  t59_g186 : AOI21D0BWP7T port map(A1 => t59_n_4, A2 => t59_n_5, B => reset, ZN => t59_n_7);
  t59_g187 : AOI22D0BWP7T port map(A1 => t59_state(1), A2 => t59_n_5, B1 => t59_state(0), B2 => t59_n_3, ZN => t59_n_6);
  t59_g188 : ND3D0BWP7T port map(A1 => yo5, A2 => xo3, A3 => t59_n_2, ZN => t59_n_5);
  t59_g189 : ND2D1BWP7T port map(A1 => t59_state(0), A2 => t59_n_2, ZN => t59_n_4);
  t59_drc_bufs : INVD0BWP7T port map(I => t59_n_3, ZN => t59_n_2);
  t59_drc_bufs192 : INVD0BWP7T port map(I => lethal, ZN => t59_n_3);
  t59_state_reg_0 : DFD1BWP7T port map(CP => clk, D => t59_n_7, Q => t59_state(0), QN => t59_n_11);
  t59_state_reg_1 : DFD1BWP7T port map(CP => clk, D => t59_n_8, Q => t59_state(1), QN => t59_n_9);
  t60_g68 : INVD4BWP7T port map(I => t60_state, ZN => y5(12));
  t60_state_reg : DFQD1BWP7T port map(CP => clk, D => t60_n_3, Q => t60_state);
  t60_g118 : AOI211XD0BWP7T port map(A1 => y5(12), A2 => t60_n_2, B => n_126, C => t60_n_1, ZN => t60_n_3);
  t60_g119 : ND2D0BWP7T port map(A1 => yo5, A2 => xo4, ZN => t60_n_2);
  t60_g120 : INVD0BWP7T port map(I => lethal, ZN => t60_n_1);
  tie_0_cell : TIELBWP7T port map(ZN => y1(19));
  tie_1_cell : TIEHBWP7T port map(Z => y0(21));

end synthesised;
