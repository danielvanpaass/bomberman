library IEEE;
use IEEE.std_logic_1164.ALL;

entity vga_top_lvl_tb is
end vga_top_lvl_tb;

