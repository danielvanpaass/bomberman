configuration playground_tb_behaviour_cfg of playground_tb is
   for behaviour
      for all: playground use configuration work.playground_behaviour_cfg;
      end for;
   end for;
end playground_tb_behaviour_cfg;
