configuration bombcook_tb_behaviour_cfg of bombcook_tb is
   for behaviour
      for all: bombcook use configuration work.bombcook_behaviour_cfg;
      end for;
   end for;
end bombcook_tb_behaviour_cfg;
