library IEEE;
use IEEE.std_logic_1164.ALL;

entity tile_fsm_crate is
   port(lethalx : in  std_logic);
end tile_fsm_crate;

