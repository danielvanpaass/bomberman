configuration hitscan_behaviour_cfg of hitscan is
   for behaviour
   end for;
end hitscan_behaviour_cfg;
