library IEEE;
use IEEE.std_logic_1164.ALL;

entity hitbox_top_lvl_tb is
end hitbox_top_lvl_tb;

