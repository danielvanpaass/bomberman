configuration tile_stdcrate_behaviour_cfg of tile_stdcrate is
   for behaviour
   end for;
end tile_stdcrate_behaviour_cfg;
