configuration reg_behaviour_cfg of reg is
   for behaviour
   end for;
end reg_behaviour_cfg;
