library IEEE;
use IEEE.std_logic_1164.ALL;

entity map_gen is
   port(crates_vector : out std_logic_vector(64 downto 0));
end map_gen;


