configuration xy_convert_behaviour_cfg of xy_convert is
   for behaviour
   end for;
end xy_convert_behaviour_cfg;
