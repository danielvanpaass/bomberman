configuration xy_convert_tb_behaviour_cfg of xy_convert_tb is
   for behaviour
      for all: xy_convert use configuration work.xy_convert_behaviour_cfg;
      end for;
   end for;
end xy_convert_tb_behaviour_cfg;
