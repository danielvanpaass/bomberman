library IEEE;
use IEEE.std_logic_1164.ALL;

architecture behaviour of sprites_tb is
   component sprites
      port(victory : in std_logic;
   playground: in  std_logic_vector(241 downto 0);
   	clk : in std_logic;
   	reset: in std_logic;
           x_p1          : in  std_logic_vector(3 downto 0);
           y_p1          : in  std_logic_vector(3 downto 0);
          x_p2          : in  std_logic_vector(3 downto 0);
          y_p2          : in  std_logic_vector(3 downto 0);
           x_bomb_a      : in  std_logic_vector(3 downto 0);
           y_bomb_a      : in  std_logic_vector(3 downto 0);
           bomb_a_enable : in  std_logic;
           x_bomb_b      : in  std_logic_vector(3 downto 0);
           y_bomb_b      : in  std_logic_vector(3 downto 0);
           bomb_b_enable : in  std_logic;
           x_bomb_c      : in  std_logic_vector(3 downto 0);
           y_bomb_c      : in  std_logic_vector(3 downto 0);
           bomb_c_enable : in  std_logic;
           x_bomb_d      : in  std_logic_vector(3 downto 0);
           y_bomb_d      : in  std_logic_vector(3 downto 0);
           bomb_d_enable : in  std_logic;
           x_bomb_e      : in  std_logic_vector(3 downto 0);
           y_bomb_e      : in  std_logic_vector(3 downto 0);
           bomb_e_enable : in  std_logic;
           x_bomb_f      : in  std_logic_vector(3 downto 0);
           y_bomb_f      : in  std_logic_vector(3 downto 0);
           bomb_f_enable : in  std_logic;
           x_bomb_g      : in  std_logic_vector(3 downto 0);
           y_bomb_g      : in  std_logic_vector(3 downto 0);
           bomb_g_enable : in  std_logic;
           x_bomb_h      : in  std_logic_vector(3 downto 0);
           y_bomb_h      : in  std_logic_vector(3 downto 0);
           bomb_h_enable : in  std_logic;
           x_map         : in  std_logic_vector(3 downto 0);
           y_map         : in  std_logic_vector(3 downto 0);
           input_h_map         : in  std_logic_vector(5 downto 0);
           input_v_map         : in  std_logic_vector(6 downto 0);
   	red : out std_logic;
   	green : out std_logic;
   	blue: out std_logic);      
   end component;
   signal victory : std_logic;
   signal playground: std_logic_vector(241 downto 0);
   signal clk : std_logic;
   signal reset: std_logic;
   signal x_p1          : std_logic_vector(3 downto 0);
   signal y_p1          : std_logic_vector(3 downto 0);
   signal x_p2          : std_logic_vector(3 downto 0);
   signal y_p2          : std_logic_vector(3 downto 0);
   signal x_bomb_a      : std_logic_vector(3 downto 0);
   signal y_bomb_a      : std_logic_vector(3 downto 0);
   signal bomb_a_enable : std_logic;
   signal x_bomb_b      : std_logic_vector(3 downto 0);
   signal y_bomb_b      : std_logic_vector(3 downto 0);
   signal bomb_b_enable : std_logic;
   signal x_bomb_c      : std_logic_vector(3 downto 0);
   signal y_bomb_c      : std_logic_vector(3 downto 0);
   signal bomb_c_enable : std_logic;
   signal x_bomb_d      : std_logic_vector(3 downto 0);
   signal y_bomb_d      : std_logic_vector(3 downto 0);
   signal bomb_d_enable : std_logic;
   signal x_bomb_e      : std_logic_vector(3 downto 0);
   signal y_bomb_e      : std_logic_vector(3 downto 0);
   signal bomb_e_enable : std_logic;
   signal x_bomb_f      : std_logic_vector(3 downto 0);
   signal y_bomb_f      : std_logic_vector(3 downto 0);
   signal bomb_f_enable : std_logic;
   signal x_bomb_g      : std_logic_vector(3 downto 0);
   signal y_bomb_g      : std_logic_vector(3 downto 0);
   signal bomb_g_enable : std_logic;
   signal x_bomb_h      : std_logic_vector(3 downto 0);
   signal y_bomb_h      : std_logic_vector(3 downto 0);
   signal bomb_h_enable : std_logic;
   signal x_map         : std_logic_vector(3 downto 0);
   signal y_map         : std_logic_vector(3 downto 0);
   signal input_h_map         : std_logic_vector(5 downto 0);
   signal input_v_map         : std_logic_vector(6 downto 0);
   signal red : std_logic;
   signal green : std_logic;
   signal blue: std_logic;
begin
test: sprites port map (victory, playground, clk, reset, x_p1, y_p1, x_p2, y_p2, x_bomb_a, y_bomb_a, bomb_a_enable, x_bomb_b, y_bomb_b, bomb_b_enable, x_bomb_c, y_bomb_c, bomb_c_enable, x_bomb_d, y_bomb_d, bomb_d_enable, x_bomb_e, y_bomb_e, bomb_e_enable, x_bomb_f, y_bomb_f, bomb_f_enable, x_bomb_g, y_bomb_g, bomb_g_enable, x_bomb_h, y_bomb_h, bomb_h_enable, x_map, y_map, input_h_map, input_v_map, red, green, blue);
   clk <= '0' after 1 ns when clk /= '0' else '1' after 1 ns;
   reset <= '1' after 0 ns,
'0' after 3 ns;   
victory <= '0' after 0 ns;
   playground(0) <= '1' after 0 ns;
   playground(1) <= '1' after 0 ns;
   playground(2) <= '1' after 0 ns;
   playground(3) <= '1' after 0 ns;
   playground(4) <= '1' after 0 ns;
   playground(5) <= '1' after 0 ns;
   playground(6) <= '1' after 0 ns;
   playground(7) <= '1' after 0 ns;
   playground(8) <= '1' after 0 ns;
   playground(9) <= '1' after 0 ns;
   playground(10) <= '1' after 0 ns;
   playground(11) <= '1' after 0 ns;
   playground(12) <= '1' after 0 ns;
   playground(13) <= '1' after 0 ns;
   playground(14) <= '1' after 0 ns;
   playground(15) <= '1' after 0 ns;
   playground(16) <= '1' after 0 ns;
   playground(17) <= '1' after 0 ns;
   playground(18) <= '1' after 0 ns;
   playground(19) <= '1' after 0 ns;
   playground(20) <= '1' after 0 ns;
   playground(21) <= '1' after 0 ns;
   playground(22) <= '1' after 0 ns;
   playground(23) <= '1' after 0 ns;
   playground(24) <= '1' after 0 ns;
   playground(25) <= '0' after 0 ns;
   playground(26) <= '1' after 0 ns;
   playground(27) <= '0' after 0 ns;
   playground(28) <= '1' after 0 ns;
   playground(29) <= '0' after 0 ns;
   playground(30) <= '1' after 0 ns;
   playground(31) <= '0' after 0 ns;
   playground(32) <= '1' after 0 ns;
   playground(33) <= '0' after 0 ns;
   playground(34) <= '1' after 0 ns;
   playground(35) <= '0' after 0 ns;
   playground(36) <= '1' after 0 ns;
   playground(37) <= '0' after 0 ns;
   playground(38) <= '1' after 0 ns;
   playground(39) <= '0' after 0 ns;
   playground(40) <= '1' after 0 ns;
   playground(41) <= '0' after 0 ns;
   playground(42) <= '1' after 0 ns;
   playground(43) <= '0' after 0 ns;
   playground(44) <= '1' after 0 ns;
   playground(45) <= '0' after 0 ns;
   playground(46) <= '0' after 0 ns;
   playground(47) <= '0' after 0 ns;
   playground(48) <= '0' after 0 ns;
   playground(49) <= '0' after 0 ns;
   playground(50) <= '0' after 0 ns;
   playground(51) <= '0' after 0 ns;
   playground(52) <= '0' after 0 ns;
   playground(53) <= '0' after 0 ns;
   playground(54) <= '0' after 0 ns;
   playground(55) <= '0' after 0 ns;
   playground(56) <= '0' after 0 ns;
   playground(57) <= '0' after 0 ns;
   playground(58) <= '0' after 0 ns;
   playground(59) <= '0' after 0 ns;
   playground(60) <= '0' after 0 ns;
   playground(61) <= '0' after 0 ns;
   playground(62) <= '0' after 0 ns;
   playground(63) <= '0' after 0 ns;
   playground(64) <= '0' after 0 ns;
   playground(65) <= '0' after 0 ns;
   playground(66) <= '0' after 0 ns;
   playground(67) <= '0' after 0 ns;
   playground(68) <= '1' after 0 ns;
   playground(69) <= '0' after 0 ns;
   playground(70) <= '1' after 0 ns;
   playground(71) <= '0' after 0 ns;
   playground(72) <= '1' after 0 ns;
   playground(73) <= '0' after 0 ns;
   playground(74) <= '1' after 0 ns;
   playground(75) <= '0' after 0 ns;
   playground(76) <= '1' after 0 ns;
   playground(77) <= '0' after 0 ns;
   playground(78) <= '1' after 0 ns;
   playground(79) <= '0' after 0 ns;
   playground(80) <= '1' after 0 ns;
   playground(81) <= '0' after 0 ns;
   playground(82) <= '1' after 0 ns;
   playground(83) <= '0' after 0 ns;
   playground(84) <= '1' after 0 ns;
   playground(85) <= '0' after 0 ns;
   playground(86) <= '1' after 0 ns;
   playground(87) <= '0' after 0 ns;
   playground(88) <= '1' after 0 ns;
   playground(89) <= '0' after 0 ns;
   playground(90) <= '0' after 0 ns;
   playground(91) <= '0' after 0 ns;
   playground(92) <= '0' after 0 ns;
   playground(93) <= '0' after 0 ns;
   playground(94) <= '0' after 0 ns;
   playground(95) <= '0' after 0 ns;
   playground(96) <= '0' after 0 ns;
   playground(97) <= '0' after 0 ns;
   playground(98) <= '0' after 0 ns;
   playground(99) <= '0' after 0 ns;
   playground(100) <= '0' after 0 ns;
   playground(101) <= '0' after 0 ns;
   playground(102) <= '0' after 0 ns;
   playground(103) <= '0' after 0 ns;
   playground(104) <= '0' after 0 ns;
   playground(105) <= '0' after 0 ns;
   playground(106) <= '0' after 0 ns;
   playground(107) <= '0' after 0 ns;
   playground(108) <= '0' after 0 ns;
   playground(109) <= '0' after 0 ns;
   playground(110) <= '0' after 0 ns;
   playground(111) <= '0' after 0 ns;
   playground(112) <= '0' after 0 ns;
   playground(113) <= '0' after 0 ns;
   playground(114) <= '0' after 0 ns;
   playground(115) <= '0' after 0 ns;
   playground(116) <= '0' after 0 ns;
   playground(117) <= '0' after 0 ns;
   playground(118) <= '0' after 0 ns;
   playground(119) <= '0' after 0 ns;
   playground(120) <= '0' after 0 ns;
   playground(121) <= '0' after 0 ns;
   playground(122) <= '0' after 0 ns;
   playground(123) <= '0' after 0 ns;
   playground(124) <= '0' after 0 ns;
   playground(125) <= '0' after 0 ns;
   playground(126) <= '0' after 0 ns;
   playground(127) <= '0' after 0 ns;
   playground(128) <= '0' after 0 ns;
   playground(129) <= '0' after 0 ns;
   playground(130) <= '0' after 0 ns;
   playground(131) <= '0' after 0 ns;
   playground(132) <= '0' after 0 ns;
   playground(133) <= '0' after 0 ns;
   playground(134) <= '0' after 0 ns;
   playground(135) <= '0' after 0 ns;
   playground(136) <= '0' after 0 ns;
   playground(137) <= '0' after 0 ns;
   playground(138) <= '0' after 0 ns;
   playground(139) <= '0' after 0 ns;
   playground(140) <= '0' after 0 ns;
   playground(141) <= '0' after 0 ns;
   playground(142) <= '0' after 0 ns;
   playground(143) <= '0' after 0 ns;
   playground(144) <= '0' after 0 ns;
   playground(145) <= '0' after 0 ns;
   playground(146) <= '0' after 0 ns;
   playground(147) <= '0' after 0 ns;
   playground(148) <= '0' after 0 ns;
   playground(149) <= '0' after 0 ns;
   playground(150) <= '0' after 0 ns;
   playground(151) <= '0' after 0 ns;
   playground(152) <= '0' after 0 ns;
   playground(153) <= '0' after 0 ns;
   playground(154) <= '0' after 0 ns;
   playground(155) <= '0' after 0 ns;
   playground(156) <= '0' after 0 ns;
   playground(157) <= '0' after 0 ns;
   playground(158) <= '0' after 0 ns;
   playground(159) <= '0' after 0 ns;
   playground(160) <= '0' after 0 ns;
   playground(161) <= '0' after 0 ns;
   playground(162) <= '0' after 0 ns;
   playground(163) <= '0' after 0 ns;
   playground(164) <= '0' after 0 ns;
   playground(165) <= '0' after 0 ns;
   playground(166) <= '0' after 0 ns;
   playground(167) <= '0' after 0 ns;
   playground(168) <= '0' after 0 ns;
   playground(169) <= '0' after 0 ns;
   playground(170) <= '0' after 0 ns;
   playground(171) <= '0' after 0 ns;
   playground(172) <= '0' after 0 ns;
   playground(173) <= '0' after 0 ns;
   playground(174) <= '0' after 0 ns;
   playground(175) <= '0' after 0 ns;
   playground(176) <= '0' after 0 ns;
   playground(177) <= '0' after 0 ns;
   playground(178) <= '0' after 0 ns;
   playground(179) <= '0' after 0 ns;
   playground(180) <= '0' after 0 ns;
   playground(181) <= '0' after 0 ns;
   playground(182) <= '0' after 0 ns;
   playground(183) <= '0' after 0 ns;
   playground(184) <= '0' after 0 ns;
   playground(185) <= '0' after 0 ns;
   playground(186) <= '0' after 0 ns;
   playground(187) <= '0' after 0 ns;
   playground(188) <= '0' after 0 ns;
   playground(189) <= '0' after 0 ns;
   playground(190) <= '0' after 0 ns;
   playground(191) <= '0' after 0 ns;
   playground(192) <= '0' after 0 ns;
   playground(193) <= '0' after 0 ns;
   playground(194) <= '0' after 0 ns;
   playground(195) <= '0' after 0 ns;
   playground(196) <= '0' after 0 ns;
   playground(197) <= '0' after 0 ns;
   playground(198) <= '0' after 0 ns;
   playground(199) <= '0' after 0 ns;
   playground(200) <= '0' after 0 ns;
   playground(201) <= '0' after 0 ns;
   playground(202) <= '0' after 0 ns;
   playground(203) <= '0' after 0 ns;
   playground(204) <= '0' after 0 ns;
   playground(205) <= '0' after 0 ns;
   playground(206) <= '0' after 0 ns;
   playground(207) <= '0' after 0 ns;
   playground(208) <= '0' after 0 ns;
   playground(209) <= '0' after 0 ns;
   playground(210) <= '0' after 0 ns;
   playground(211) <= '0' after 0 ns;
   playground(212) <= '0' after 0 ns;
   playground(213) <= '0' after 0 ns;
   playground(214) <= '0' after 0 ns;
   playground(215) <= '0' after 0 ns;
   playground(216) <= '0' after 0 ns;
   playground(217) <= '0' after 0 ns;
   playground(218) <= '0' after 0 ns;
   playground(219) <= '0' after 0 ns;
   playground(220) <= '1' after 0 ns;
   playground(221) <= '1' after 0 ns;
   playground(222) <= '1' after 0 ns;
   playground(223) <= '1' after 0 ns;
   playground(224) <= '1' after 0 ns;
   playground(225) <= '1' after 0 ns;
   playground(226) <= '1' after 0 ns;
   playground(227) <= '1' after 0 ns;
   playground(228) <= '1' after 0 ns;
   playground(229) <= '1' after 0 ns;
   playground(230) <= '1' after 0 ns;
   playground(231) <= '1' after 0 ns;
   playground(232) <= '1' after 0 ns;
   playground(233) <= '1' after 0 ns;
   playground(234) <= '1' after 0 ns;
   playground(235) <= '1' after 0 ns;
   playground(236) <= '1' after 0 ns;
   playground(237) <= '1' after 0 ns;
   playground(238) <= '1' after 0 ns;
   playground(239) <= '1' after 0 ns;
   playground(240) <= '0' after 0 ns;
   playground(241) <= '0' after 0 ns;
   x_p1(0) <= '0' after 0 ns;
   x_p1(1) <= '0' after 0 ns;
   x_p1(2) <= '0' after 0 ns;
   x_p1(3) <= '0' after 0 ns;
   y_p1(0) <= '0' after 0 ns;
   y_p1(1) <= '0' after 0 ns;
   y_p1(2) <= '0' after 0 ns;
   y_p1(3) <= '0' after 0 ns;
   x_p2(0) <= '1' after 0 ns;
   x_p2(1) <= '1' after 0 ns;
   x_p2(2) <= '1' after 0 ns;
   x_p2(3) <= '1' after 0 ns;
   y_p2(0) <= '1' after 0 ns;
   y_p2(1) <= '1' after 0 ns;
   y_p2(2) <= '1' after 0 ns;
   y_p2(3) <= '1' after 0 ns;
   x_bomb_a(0) <= '0' after 0 ns;
   x_bomb_a(1) <= '0' after 0 ns;
   x_bomb_a(2) <= '0' after 0 ns;
   x_bomb_a(3) <= '0' after 0 ns;
   y_bomb_a(0) <= '0' after 0 ns;
   y_bomb_a(1) <= '0' after 0 ns;
   y_bomb_a(2) <= '0' after 0 ns;
   y_bomb_a(3) <= '0' after 0 ns;
   bomb_a_enable <= '1' after 0 ns;
   x_bomb_b(0) <= '0' after 0 ns;
   x_bomb_b(1) <= '0' after 0 ns;
   x_bomb_b(2) <= '0' after 0 ns;
   x_bomb_b(3) <= '0' after 0 ns;
   y_bomb_b(0) <= '0' after 0 ns;
   y_bomb_b(1) <= '0' after 0 ns;
   y_bomb_b(2) <= '0' after 0 ns;
   y_bomb_b(3) <= '0' after 0 ns;
   bomb_b_enable <= '0' after 0 ns;
   x_bomb_c(0) <= '0' after 0 ns;
   x_bomb_c(1) <= '0' after 0 ns;
   x_bomb_c(2) <= '0' after 0 ns;
   x_bomb_c(3) <= '0' after 0 ns;
   y_bomb_c(0) <= '0' after 0 ns;
   y_bomb_c(1) <= '0' after 0 ns;
   y_bomb_c(2) <= '0' after 0 ns;
   y_bomb_c(3) <= '0' after 0 ns;
   bomb_c_enable <= '0' after 0 ns;
   x_bomb_d(0) <= '0' after 0 ns;
   x_bomb_d(1) <= '0' after 0 ns;
   x_bomb_d(2) <= '0' after 0 ns;
   x_bomb_d(3) <= '0' after 0 ns;
   y_bomb_d(0) <= '0' after 0 ns;
   y_bomb_d(1) <= '0' after 0 ns;
   y_bomb_d(2) <= '0' after 0 ns;
   y_bomb_d(3) <= '0' after 0 ns;
   bomb_d_enable <= '0' after 0 ns;
   x_bomb_e(0) <= '0' after 0 ns;
   x_bomb_e(1) <= '0' after 0 ns;
   x_bomb_e(2) <= '0' after 0 ns;
   x_bomb_e(3) <= '0' after 0 ns;
   y_bomb_e(0) <= '0' after 0 ns;
   y_bomb_e(1) <= '0' after 0 ns;
   y_bomb_e(2) <= '0' after 0 ns;
   y_bomb_e(3) <= '0' after 0 ns;
   bomb_e_enable <= '0' after 0 ns;
   x_bomb_f(0) <= '0' after 0 ns;
   x_bomb_f(1) <= '0' after 0 ns;
   x_bomb_f(2) <= '0' after 0 ns;
   x_bomb_f(3) <= '0' after 0 ns;
   y_bomb_f(0) <= '0' after 0 ns;
   y_bomb_f(1) <= '0' after 0 ns;
   y_bomb_f(2) <= '0' after 0 ns;
   y_bomb_f(3) <= '0' after 0 ns;
   bomb_f_enable <= '0' after 0 ns;
   x_bomb_g(0) <= '0' after 0 ns;
   x_bomb_g(1) <= '0' after 0 ns;
   x_bomb_g(2) <= '0' after 0 ns;
   x_bomb_g(3) <= '0' after 0 ns;
   y_bomb_g(0) <= '0' after 0 ns;
   y_bomb_g(1) <= '0' after 0 ns;
   y_bomb_g(2) <= '0' after 0 ns;
   y_bomb_g(3) <= '0' after 0 ns;
   bomb_g_enable <= '0' after 0 ns;
   x_bomb_h(0) <= '0' after 0 ns;
   x_bomb_h(1) <= '0' after 0 ns;
   x_bomb_h(2) <= '0' after 0 ns;
   x_bomb_h(3) <= '0' after 0 ns;
   y_bomb_h(0) <= '0' after 0 ns;
   y_bomb_h(1) <= '0' after 0 ns;
   y_bomb_h(2) <= '0' after 0 ns;
   y_bomb_h(3) <= '0' after 0 ns;
   bomb_h_enable <= '0' after 0 ns;
   x_map <= "0000" after 0 ns;
   y_map <= "0000" after 0 ns;
	--"0001" after 9600 ns,
	--"0010" after 19200 ns;

   y_map(1) <= '0' after 0 ns;
   y_map(2) <= '0' after 0 ns;
   y_map(3) <= '0' after 0 ns;
  input_h_map(0) <= '0' after 0 ns,
      '1' after 10 ns when  input_h_map(0)/= '1' else '0' after 10 ns;

   input_h_map(1) <= '0' after 0 ns,
      '1' after 20 ns when input_h_map(1) /= '1' else '0' after 20 ns;

   input_h_map(2) <= '0' after 0 ns,
      '1' after 40 ns when input_h_map(2) /= '1' else '0' after 40 ns;

   input_h_map(3) <= '0' after 0 ns,
      '1' after 80 ns when input_h_map(3) /= '1' else '0' after 80 ns;

   input_h_map(4) <= '0' after 0 ns,
      '1' after 160 ns when input_h_map(4) /= '1' else '0' after 160 ns;

   input_h_map(5) <= '0' after 0 ns;

   input_v_map(0) <= '0' after 0 ns,
      '1' after 320 ns when input_v_map(0) /= '1' else '0' after 320 ns;

   input_v_map(1) <= '0' after 0 ns,
	'1' after 640 ns when input_v_map(1) /= '1' else '0' after 640 ns;

   input_v_map(2) <= '0' after 0 ns,
	'1' after 1280 ns when input_v_map(2) /= '1' else '0' after 1280 ns;

   input_v_map(3) <= '0' after 0 ns,
	'1' after 2560 ns when input_v_map(3) /= '1' else '0' after 2560 ns;

   input_v_map(4) <= '0' after 0 ns,
	'1' after 5120 ns when input_v_map(4) /= '1' else '0' after 5120 ns;

   input_v_map(5) <= '0' after 0 ns,
	'1' after 10240 ns when input_v_map(5) /= '1' else '0' after 10240 ns; 

    input_v_map(6)<= '0' after 0 ns;
end behaviour;
