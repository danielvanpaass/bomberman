configuration ff2_behaviour_cfg of ff2 is
   for behaviour
   end for;
end ff2_behaviour_cfg;
