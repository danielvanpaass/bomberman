configuration playground_behaviour_cfg of playground is
   for behaviour
      for all: tile_stdempty use configuration work.tile_stdempty_behaviour_cfg;
      end for;
   end for;
end playground_behaviour_cfg;
