library IEEE;
use IEEE.std_logic_1164.ALL;

entity bombcook_tb is
end bombcook_tb;

