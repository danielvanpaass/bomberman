library IEEE;
use IEEE.std_logic_1164.ALL;

entity playground_tb is
end playground_tb;

