configuration selector_behaviour_cfg of selector is
   for behaviour
   end for;
end selector_behaviour_cfg;
