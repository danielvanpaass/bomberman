configuration hitbox_tb_behaviour_directions_cfg of hitbox_tb is
   for behaviour_directions
      for all: hitbox use configuration work.hitbox_hitbox_behaviour_cfg;
      end for;
   end for;
end hitbox_tb_behaviour_directions_cfg;
