
library ieee;
use ieee.std_logic_1164.all;
--library tcb018gbwp7t;
--use tcb018gbwp7t.all;

architecture synthesised of obstacle_map is

  component BUFFD4BWP7T
    port(I : in std_logic; Z : out std_logic);
  end component;


begin

  drc_bufs : BUFFD4BWP7T port map(I => playground(221), Z => obstacle(110));
  drc_bufs3 : BUFFD4BWP7T port map(I => playground(21), Z => obstacle(10));
  drc_bufs6 : BUFFD4BWP7T port map(I => playground(19), Z => obstacle(9));
  drc_bufs9 : BUFFD4BWP7T port map(I => playground(17), Z => obstacle(8));
  drc_bufs12 : BUFFD4BWP7T port map(I => playground(15), Z => obstacle(7));
  drc_bufs15 : BUFFD4BWP7T port map(I => playground(13), Z => obstacle(6));
  drc_bufs18 : BUFFD4BWP7T port map(I => playground(11), Z => obstacle(5));
  drc_bufs21 : BUFFD4BWP7T port map(I => playground(9), Z => obstacle(4));
  drc_bufs24 : BUFFD4BWP7T port map(I => playground(7), Z => obstacle(3));
  drc_bufs27 : BUFFD4BWP7T port map(I => playground(5), Z => obstacle(2));
  drc_bufs30 : BUFFD4BWP7T port map(I => playground(3), Z => obstacle(1));
  drc_bufs33 : BUFFD4BWP7T port map(I => playground(1), Z => obstacle(0));
  drc_bufs36 : BUFFD4BWP7T port map(I => playground(43), Z => obstacle(21));
  drc_bufs39 : BUFFD4BWP7T port map(I => playground(41), Z => obstacle(20));
  drc_bufs42 : BUFFD4BWP7T port map(I => playground(39), Z => obstacle(19));
  drc_bufs45 : BUFFD4BWP7T port map(I => playground(37), Z => obstacle(18));
  drc_bufs48 : BUFFD4BWP7T port map(I => playground(35), Z => obstacle(17));
  drc_bufs51 : BUFFD4BWP7T port map(I => playground(33), Z => obstacle(16));
  drc_bufs54 : BUFFD4BWP7T port map(I => playground(31), Z => obstacle(15));
  drc_bufs57 : BUFFD4BWP7T port map(I => playground(29), Z => obstacle(14));
  drc_bufs60 : BUFFD4BWP7T port map(I => playground(27), Z => obstacle(13));
  drc_bufs63 : BUFFD4BWP7T port map(I => playground(25), Z => obstacle(12));
  drc_bufs66 : BUFFD4BWP7T port map(I => playground(23), Z => obstacle(11));
  drc_bufs69 : BUFFD4BWP7T port map(I => playground(65), Z => obstacle(32));
  drc_bufs72 : BUFFD4BWP7T port map(I => playground(63), Z => obstacle(31));
  drc_bufs75 : BUFFD4BWP7T port map(I => playground(61), Z => obstacle(30));
  drc_bufs78 : BUFFD4BWP7T port map(I => playground(59), Z => obstacle(29));
  drc_bufs81 : BUFFD4BWP7T port map(I => playground(57), Z => obstacle(28));
  drc_bufs84 : BUFFD4BWP7T port map(I => playground(55), Z => obstacle(27));
  drc_bufs87 : BUFFD4BWP7T port map(I => playground(53), Z => obstacle(26));
  drc_bufs90 : BUFFD4BWP7T port map(I => playground(51), Z => obstacle(25));
  drc_bufs93 : BUFFD4BWP7T port map(I => playground(49), Z => obstacle(24));
  drc_bufs96 : BUFFD4BWP7T port map(I => playground(47), Z => obstacle(23));
  drc_bufs99 : BUFFD4BWP7T port map(I => playground(45), Z => obstacle(22));
  drc_bufs102 : BUFFD4BWP7T port map(I => playground(87), Z => obstacle(43));
  drc_bufs105 : BUFFD4BWP7T port map(I => playground(85), Z => obstacle(42));
  drc_bufs108 : BUFFD4BWP7T port map(I => playground(83), Z => obstacle(41));
  drc_bufs111 : BUFFD4BWP7T port map(I => playground(81), Z => obstacle(40));
  drc_bufs114 : BUFFD4BWP7T port map(I => playground(79), Z => obstacle(39));
  drc_bufs117 : BUFFD4BWP7T port map(I => playground(77), Z => obstacle(38));
  drc_bufs120 : BUFFD4BWP7T port map(I => playground(75), Z => obstacle(37));
  drc_bufs123 : BUFFD4BWP7T port map(I => playground(73), Z => obstacle(36));
  drc_bufs126 : BUFFD4BWP7T port map(I => playground(71), Z => obstacle(35));
  drc_bufs129 : BUFFD4BWP7T port map(I => playground(69), Z => obstacle(34));
  drc_bufs132 : BUFFD4BWP7T port map(I => playground(67), Z => obstacle(33));
  drc_bufs135 : BUFFD4BWP7T port map(I => playground(109), Z => obstacle(54));
  drc_bufs138 : BUFFD4BWP7T port map(I => playground(107), Z => obstacle(53));
  drc_bufs141 : BUFFD4BWP7T port map(I => playground(105), Z => obstacle(52));
  drc_bufs144 : BUFFD4BWP7T port map(I => playground(103), Z => obstacle(51));
  drc_bufs147 : BUFFD4BWP7T port map(I => playground(101), Z => obstacle(50));
  drc_bufs150 : BUFFD4BWP7T port map(I => playground(99), Z => obstacle(49));
  drc_bufs153 : BUFFD4BWP7T port map(I => playground(97), Z => obstacle(48));
  drc_bufs156 : BUFFD4BWP7T port map(I => playground(95), Z => obstacle(47));
  drc_bufs159 : BUFFD4BWP7T port map(I => playground(93), Z => obstacle(46));
  drc_bufs162 : BUFFD4BWP7T port map(I => playground(91), Z => obstacle(45));
  drc_bufs165 : BUFFD4BWP7T port map(I => playground(89), Z => obstacle(44));
  drc_bufs168 : BUFFD4BWP7T port map(I => playground(131), Z => obstacle(65));
  drc_bufs171 : BUFFD4BWP7T port map(I => playground(129), Z => obstacle(64));
  drc_bufs174 : BUFFD4BWP7T port map(I => playground(127), Z => obstacle(63));
  drc_bufs177 : BUFFD4BWP7T port map(I => playground(125), Z => obstacle(62));
  drc_bufs180 : BUFFD4BWP7T port map(I => playground(123), Z => obstacle(61));
  drc_bufs183 : BUFFD4BWP7T port map(I => playground(121), Z => obstacle(60));
  drc_bufs186 : BUFFD4BWP7T port map(I => playground(119), Z => obstacle(59));
  drc_bufs189 : BUFFD4BWP7T port map(I => playground(117), Z => obstacle(58));
  drc_bufs192 : BUFFD4BWP7T port map(I => playground(115), Z => obstacle(57));
  drc_bufs195 : BUFFD4BWP7T port map(I => playground(113), Z => obstacle(56));
  drc_bufs198 : BUFFD4BWP7T port map(I => playground(111), Z => obstacle(55));
  drc_bufs201 : BUFFD4BWP7T port map(I => playground(153), Z => obstacle(76));
  drc_bufs204 : BUFFD4BWP7T port map(I => playground(151), Z => obstacle(75));
  drc_bufs207 : BUFFD4BWP7T port map(I => playground(149), Z => obstacle(74));
  drc_bufs210 : BUFFD4BWP7T port map(I => playground(147), Z => obstacle(73));
  drc_bufs213 : BUFFD4BWP7T port map(I => playground(145), Z => obstacle(72));
  drc_bufs216 : BUFFD4BWP7T port map(I => playground(143), Z => obstacle(71));
  drc_bufs219 : BUFFD4BWP7T port map(I => playground(141), Z => obstacle(70));
  drc_bufs222 : BUFFD4BWP7T port map(I => playground(139), Z => obstacle(69));
  drc_bufs225 : BUFFD4BWP7T port map(I => playground(137), Z => obstacle(68));
  drc_bufs228 : BUFFD4BWP7T port map(I => playground(135), Z => obstacle(67));
  drc_bufs231 : BUFFD4BWP7T port map(I => playground(133), Z => obstacle(66));
  drc_bufs234 : BUFFD4BWP7T port map(I => playground(175), Z => obstacle(87));
  drc_bufs237 : BUFFD4BWP7T port map(I => playground(173), Z => obstacle(86));
  drc_bufs240 : BUFFD4BWP7T port map(I => playground(171), Z => obstacle(85));
  drc_bufs243 : BUFFD4BWP7T port map(I => playground(169), Z => obstacle(84));
  drc_bufs246 : BUFFD4BWP7T port map(I => playground(167), Z => obstacle(83));
  drc_bufs249 : BUFFD4BWP7T port map(I => playground(165), Z => obstacle(82));
  drc_bufs252 : BUFFD4BWP7T port map(I => playground(163), Z => obstacle(81));
  drc_bufs255 : BUFFD4BWP7T port map(I => playground(161), Z => obstacle(80));
  drc_bufs258 : BUFFD4BWP7T port map(I => playground(159), Z => obstacle(79));
  drc_bufs261 : BUFFD4BWP7T port map(I => playground(157), Z => obstacle(78));
  drc_bufs264 : BUFFD4BWP7T port map(I => playground(155), Z => obstacle(77));
  drc_bufs267 : BUFFD4BWP7T port map(I => playground(197), Z => obstacle(98));
  drc_bufs270 : BUFFD4BWP7T port map(I => playground(195), Z => obstacle(97));
  drc_bufs273 : BUFFD4BWP7T port map(I => playground(193), Z => obstacle(96));
  drc_bufs276 : BUFFD4BWP7T port map(I => playground(191), Z => obstacle(95));
  drc_bufs279 : BUFFD4BWP7T port map(I => playground(189), Z => obstacle(94));
  drc_bufs282 : BUFFD4BWP7T port map(I => playground(187), Z => obstacle(93));
  drc_bufs285 : BUFFD4BWP7T port map(I => playground(185), Z => obstacle(92));
  drc_bufs288 : BUFFD4BWP7T port map(I => playground(183), Z => obstacle(91));
  drc_bufs291 : BUFFD4BWP7T port map(I => playground(181), Z => obstacle(90));
  drc_bufs294 : BUFFD4BWP7T port map(I => playground(179), Z => obstacle(89));
  drc_bufs297 : BUFFD4BWP7T port map(I => playground(177), Z => obstacle(88));
  drc_bufs300 : BUFFD4BWP7T port map(I => playground(219), Z => obstacle(109));
  drc_bufs303 : BUFFD4BWP7T port map(I => playground(217), Z => obstacle(108));
  drc_bufs306 : BUFFD4BWP7T port map(I => playground(215), Z => obstacle(107));
  drc_bufs309 : BUFFD4BWP7T port map(I => playground(213), Z => obstacle(106));
  drc_bufs312 : BUFFD4BWP7T port map(I => playground(211), Z => obstacle(105));
  drc_bufs315 : BUFFD4BWP7T port map(I => playground(209), Z => obstacle(104));
  drc_bufs318 : BUFFD4BWP7T port map(I => playground(207), Z => obstacle(103));
  drc_bufs321 : BUFFD4BWP7T port map(I => playground(205), Z => obstacle(102));
  drc_bufs324 : BUFFD4BWP7T port map(I => playground(203), Z => obstacle(101));
  drc_bufs327 : BUFFD4BWP7T port map(I => playground(201), Z => obstacle(100));
  drc_bufs330 : BUFFD4BWP7T port map(I => playground(199), Z => obstacle(99));
  drc_bufs333 : BUFFD4BWP7T port map(I => playground(241), Z => obstacle(120));
  drc_bufs336 : BUFFD4BWP7T port map(I => playground(239), Z => obstacle(119));
  drc_bufs339 : BUFFD4BWP7T port map(I => playground(237), Z => obstacle(118));
  drc_bufs342 : BUFFD4BWP7T port map(I => playground(235), Z => obstacle(117));
  drc_bufs345 : BUFFD4BWP7T port map(I => playground(233), Z => obstacle(116));
  drc_bufs348 : BUFFD4BWP7T port map(I => playground(231), Z => obstacle(115));
  drc_bufs351 : BUFFD4BWP7T port map(I => playground(229), Z => obstacle(114));
  drc_bufs354 : BUFFD4BWP7T port map(I => playground(227), Z => obstacle(113));
  drc_bufs357 : BUFFD4BWP7T port map(I => playground(225), Z => obstacle(112));
  drc_bufs360 : BUFFD4BWP7T port map(I => playground(223), Z => obstacle(111));

end synthesised;
