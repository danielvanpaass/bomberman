configuration tile_stdempty_behaviour_cfg of tile_stdempty is
   for behaviour
   end for;
end tile_stdempty_behaviour_cfg;
