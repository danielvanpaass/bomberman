configuration tile_stdcrate_tb_behaviour_cfg of tile_stdcrate_tb is
   for behaviour
      for all: tile_stdcrate use configuration work.tile_stdcrate_behaviour_cfg;
      end for;
   end for;
end tile_stdcrate_tb_behaviour_cfg;
