library IEEE;
use IEEE.std_logic_1164.ALL;

entity xy_convert_tb is
end xy_convert_tb;

