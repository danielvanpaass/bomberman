configuration bomb_select_behaviour_cfg of bomb_select is
   for behaviour
   end for;
end bomb_select_behaviour_cfg;
