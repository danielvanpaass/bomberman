library IEEE;
use IEEE.std_logic_1164.ALL;

entity bomb_select_tb is
end bomb_select_tb;

